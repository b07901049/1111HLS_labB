`timescale 1 ns / 1 ps

module AESL_deadlock_detector (
    input dl_reset,
    input all_finish,
    input dl_clock);

    wire [0:0] proc_0_data_FIFO_blk;
    wire [0:0] proc_0_data_PIPO_blk;
    wire [0:0] proc_0_start_FIFO_blk;
    wire [0:0] proc_0_TLF_FIFO_blk;
    wire [0:0] proc_0_input_sync_blk;
    wire [0:0] proc_0_output_sync_blk;
    wire [0:0] proc_dep_vld_vec_0;
    reg [0:0] proc_dep_vld_vec_0_reg;
    wire [0:0] in_chan_dep_vld_vec_0;
    wire [1:0] in_chan_dep_data_vec_0;
    wire [0:0] token_in_vec_0;
    wire [0:0] out_chan_dep_vld_vec_0;
    wire [1:0] out_chan_dep_data_0;
    wire [0:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [1:0] dep_chan_data_1_0;
    wire token_1_0;
    wire [0:0] proc_1_data_FIFO_blk;
    wire [0:0] proc_1_data_PIPO_blk;
    wire [0:0] proc_1_start_FIFO_blk;
    wire [0:0] proc_1_TLF_FIFO_blk;
    wire [0:0] proc_1_input_sync_blk;
    wire [0:0] proc_1_output_sync_blk;
    wire [0:0] proc_dep_vld_vec_1;
    reg [0:0] proc_dep_vld_vec_1_reg;
    wire [0:0] in_chan_dep_vld_vec_1;
    wire [1:0] in_chan_dep_data_vec_1;
    wire [0:0] token_in_vec_1;
    wire [0:0] out_chan_dep_vld_vec_1;
    wire [1:0] out_chan_dep_data_1;
    wire [0:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [1:0] dep_chan_data_0_1;
    wire token_0_1;
    wire [1:0] dl_in_vec;
    wire dl_detect_out;
    wire token_clear;
    wire [1:0] origin;

    reg ap_done_reg_0;// for module AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            ap_done_reg_0 <= 'b0;
        end
        else begin
            ap_done_reg_0 <= AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_done & ~AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_continue;
        end
    end

    // Process: AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0
    AESL_deadlock_detect_unit #(2, 0, 1, 1) AESL_deadlock_detect_unit_0 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_0_data_FIFO_blk[0] = 1'b0;
    assign proc_0_data_PIPO_blk[0] = 1'b0;
    assign proc_0_start_FIFO_blk[0] = 1'b0;
    assign proc_0_TLF_FIFO_blk[0] = 1'b0;
    assign proc_0_input_sync_blk[0] = 1'b0 | (AESL_inst_dft.ap_sync_Loop_VITIS_LOOP_16_1_proc_U0_ap_ready & AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_idle & ~AESL_inst_dft.ap_sync_Loop_VITIS_LOOP_21_2_proc_U0_ap_ready);
    assign proc_0_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (proc_0_data_FIFO_blk[0] | proc_0_data_PIPO_blk[0] | proc_0_start_FIFO_blk[0] | proc_0_TLF_FIFO_blk[0] | proc_0_input_sync_blk[0] | proc_0_output_sync_blk[0]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[1 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[0];

    // Process: AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0
    AESL_deadlock_detect_unit #(2, 1, 1, 1) AESL_deadlock_detect_unit_1 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_1_data_FIFO_blk[0] = 1'b0;
    assign proc_1_data_PIPO_blk[0] = 1'b0;
    assign proc_1_start_FIFO_blk[0] = 1'b0;
    assign proc_1_TLF_FIFO_blk[0] = 1'b0 | (~AESL_inst_dft.temp_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_loc_channel_U.if_write) | (~AESL_inst_dft.temp_1_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_1_loc_channel_U.if_write) | (~AESL_inst_dft.temp_2_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_2_loc_channel_U.if_write) | (~AESL_inst_dft.temp_3_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_3_loc_channel_U.if_write) | (~AESL_inst_dft.temp_4_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_4_loc_channel_U.if_write) | (~AESL_inst_dft.temp_5_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_5_loc_channel_U.if_write) | (~AESL_inst_dft.temp_6_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_6_loc_channel_U.if_write) | (~AESL_inst_dft.temp_7_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_7_loc_channel_U.if_write) | (~AESL_inst_dft.temp_8_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_8_loc_channel_U.if_write) | (~AESL_inst_dft.temp_9_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_9_loc_channel_U.if_write) | (~AESL_inst_dft.temp_10_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_10_loc_channel_U.if_write) | (~AESL_inst_dft.temp_11_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_11_loc_channel_U.if_write) | (~AESL_inst_dft.temp_12_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_12_loc_channel_U.if_write) | (~AESL_inst_dft.temp_13_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_13_loc_channel_U.if_write) | (~AESL_inst_dft.temp_14_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_14_loc_channel_U.if_write) | (~AESL_inst_dft.temp_15_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_15_loc_channel_U.if_write) | (~AESL_inst_dft.temp_16_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_16_loc_channel_U.if_write) | (~AESL_inst_dft.temp_17_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_17_loc_channel_U.if_write) | (~AESL_inst_dft.temp_18_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_18_loc_channel_U.if_write) | (~AESL_inst_dft.temp_19_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_19_loc_channel_U.if_write) | (~AESL_inst_dft.temp_20_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_20_loc_channel_U.if_write) | (~AESL_inst_dft.temp_21_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_21_loc_channel_U.if_write) | (~AESL_inst_dft.temp_22_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_22_loc_channel_U.if_write) | (~AESL_inst_dft.temp_23_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_23_loc_channel_U.if_write) | (~AESL_inst_dft.temp_24_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_24_loc_channel_U.if_write) | (~AESL_inst_dft.temp_25_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_25_loc_channel_U.if_write) | (~AESL_inst_dft.temp_26_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_26_loc_channel_U.if_write) | (~AESL_inst_dft.temp_27_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_27_loc_channel_U.if_write) | (~AESL_inst_dft.temp_28_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_28_loc_channel_U.if_write) | (~AESL_inst_dft.temp_29_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_29_loc_channel_U.if_write) | (~AESL_inst_dft.temp_30_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_30_loc_channel_U.if_write) | (~AESL_inst_dft.temp_31_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_31_loc_channel_U.if_write) | (~AESL_inst_dft.temp_32_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_32_loc_channel_U.if_write) | (~AESL_inst_dft.temp_33_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_33_loc_channel_U.if_write) | (~AESL_inst_dft.temp_34_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_34_loc_channel_U.if_write) | (~AESL_inst_dft.temp_35_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_35_loc_channel_U.if_write) | (~AESL_inst_dft.temp_36_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_36_loc_channel_U.if_write) | (~AESL_inst_dft.temp_37_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_37_loc_channel_U.if_write) | (~AESL_inst_dft.temp_38_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_38_loc_channel_U.if_write) | (~AESL_inst_dft.temp_39_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_39_loc_channel_U.if_write) | (~AESL_inst_dft.temp_40_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_40_loc_channel_U.if_write) | (~AESL_inst_dft.temp_41_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_41_loc_channel_U.if_write) | (~AESL_inst_dft.temp_42_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_42_loc_channel_U.if_write) | (~AESL_inst_dft.temp_43_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_43_loc_channel_U.if_write) | (~AESL_inst_dft.temp_44_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_44_loc_channel_U.if_write) | (~AESL_inst_dft.temp_45_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_45_loc_channel_U.if_write) | (~AESL_inst_dft.temp_46_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_46_loc_channel_U.if_write) | (~AESL_inst_dft.temp_47_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_47_loc_channel_U.if_write) | (~AESL_inst_dft.temp_48_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_48_loc_channel_U.if_write) | (~AESL_inst_dft.temp_49_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_49_loc_channel_U.if_write) | (~AESL_inst_dft.temp_50_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_50_loc_channel_U.if_write) | (~AESL_inst_dft.temp_51_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_51_loc_channel_U.if_write) | (~AESL_inst_dft.temp_52_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_52_loc_channel_U.if_write) | (~AESL_inst_dft.temp_53_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_53_loc_channel_U.if_write) | (~AESL_inst_dft.temp_54_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_54_loc_channel_U.if_write) | (~AESL_inst_dft.temp_55_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_55_loc_channel_U.if_write) | (~AESL_inst_dft.temp_56_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_56_loc_channel_U.if_write) | (~AESL_inst_dft.temp_57_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_57_loc_channel_U.if_write) | (~AESL_inst_dft.temp_58_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_58_loc_channel_U.if_write) | (~AESL_inst_dft.temp_59_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_59_loc_channel_U.if_write) | (~AESL_inst_dft.temp_60_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_60_loc_channel_U.if_write) | (~AESL_inst_dft.temp_61_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_61_loc_channel_U.if_write) | (~AESL_inst_dft.temp_62_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_62_loc_channel_U.if_write) | (~AESL_inst_dft.temp_63_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_63_loc_channel_U.if_write) | (~AESL_inst_dft.temp_64_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_64_loc_channel_U.if_write) | (~AESL_inst_dft.temp_65_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_65_loc_channel_U.if_write) | (~AESL_inst_dft.temp_66_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_66_loc_channel_U.if_write) | (~AESL_inst_dft.temp_67_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_67_loc_channel_U.if_write) | (~AESL_inst_dft.temp_68_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_68_loc_channel_U.if_write) | (~AESL_inst_dft.temp_69_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_69_loc_channel_U.if_write) | (~AESL_inst_dft.temp_70_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_70_loc_channel_U.if_write) | (~AESL_inst_dft.temp_71_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_71_loc_channel_U.if_write) | (~AESL_inst_dft.temp_72_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_72_loc_channel_U.if_write) | (~AESL_inst_dft.temp_73_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_73_loc_channel_U.if_write) | (~AESL_inst_dft.temp_74_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_74_loc_channel_U.if_write) | (~AESL_inst_dft.temp_75_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_75_loc_channel_U.if_write) | (~AESL_inst_dft.temp_76_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_76_loc_channel_U.if_write) | (~AESL_inst_dft.temp_77_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_77_loc_channel_U.if_write) | (~AESL_inst_dft.temp_78_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_78_loc_channel_U.if_write) | (~AESL_inst_dft.temp_79_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_79_loc_channel_U.if_write) | (~AESL_inst_dft.temp_80_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_80_loc_channel_U.if_write) | (~AESL_inst_dft.temp_81_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_81_loc_channel_U.if_write) | (~AESL_inst_dft.temp_82_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_82_loc_channel_U.if_write) | (~AESL_inst_dft.temp_83_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_83_loc_channel_U.if_write) | (~AESL_inst_dft.temp_84_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_84_loc_channel_U.if_write) | (~AESL_inst_dft.temp_85_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_85_loc_channel_U.if_write) | (~AESL_inst_dft.temp_86_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_86_loc_channel_U.if_write) | (~AESL_inst_dft.temp_87_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_87_loc_channel_U.if_write) | (~AESL_inst_dft.temp_88_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_88_loc_channel_U.if_write) | (~AESL_inst_dft.temp_89_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_89_loc_channel_U.if_write) | (~AESL_inst_dft.temp_90_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_90_loc_channel_U.if_write) | (~AESL_inst_dft.temp_91_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_91_loc_channel_U.if_write) | (~AESL_inst_dft.temp_92_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_92_loc_channel_U.if_write) | (~AESL_inst_dft.temp_93_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_93_loc_channel_U.if_write) | (~AESL_inst_dft.temp_94_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_94_loc_channel_U.if_write) | (~AESL_inst_dft.temp_95_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_95_loc_channel_U.if_write) | (~AESL_inst_dft.temp_96_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_96_loc_channel_U.if_write) | (~AESL_inst_dft.temp_97_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_97_loc_channel_U.if_write) | (~AESL_inst_dft.temp_98_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_98_loc_channel_U.if_write) | (~AESL_inst_dft.temp_99_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_99_loc_channel_U.if_write) | (~AESL_inst_dft.temp_100_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_100_loc_channel_U.if_write) | (~AESL_inst_dft.temp_101_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_101_loc_channel_U.if_write) | (~AESL_inst_dft.temp_102_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_102_loc_channel_U.if_write) | (~AESL_inst_dft.temp_103_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_103_loc_channel_U.if_write) | (~AESL_inst_dft.temp_104_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_104_loc_channel_U.if_write) | (~AESL_inst_dft.temp_105_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_105_loc_channel_U.if_write) | (~AESL_inst_dft.temp_106_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_106_loc_channel_U.if_write) | (~AESL_inst_dft.temp_107_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_107_loc_channel_U.if_write) | (~AESL_inst_dft.temp_108_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_108_loc_channel_U.if_write) | (~AESL_inst_dft.temp_109_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_109_loc_channel_U.if_write) | (~AESL_inst_dft.temp_110_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_110_loc_channel_U.if_write) | (~AESL_inst_dft.temp_111_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_111_loc_channel_U.if_write) | (~AESL_inst_dft.temp_112_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_112_loc_channel_U.if_write) | (~AESL_inst_dft.temp_113_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_113_loc_channel_U.if_write) | (~AESL_inst_dft.temp_114_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_114_loc_channel_U.if_write) | (~AESL_inst_dft.temp_115_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_115_loc_channel_U.if_write) | (~AESL_inst_dft.temp_116_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_116_loc_channel_U.if_write) | (~AESL_inst_dft.temp_117_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_117_loc_channel_U.if_write) | (~AESL_inst_dft.temp_118_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_118_loc_channel_U.if_write) | (~AESL_inst_dft.temp_119_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_119_loc_channel_U.if_write) | (~AESL_inst_dft.temp_120_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_120_loc_channel_U.if_write) | (~AESL_inst_dft.temp_121_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_121_loc_channel_U.if_write) | (~AESL_inst_dft.temp_122_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_122_loc_channel_U.if_write) | (~AESL_inst_dft.temp_123_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_123_loc_channel_U.if_write) | (~AESL_inst_dft.temp_124_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_124_loc_channel_U.if_write) | (~AESL_inst_dft.temp_125_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_125_loc_channel_U.if_write) | (~AESL_inst_dft.temp_126_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_126_loc_channel_U.if_write) | (~AESL_inst_dft.temp_127_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_127_loc_channel_U.if_write) | (~AESL_inst_dft.temp_128_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_128_loc_channel_U.if_write) | (~AESL_inst_dft.temp_129_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_129_loc_channel_U.if_write) | (~AESL_inst_dft.temp_130_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_130_loc_channel_U.if_write) | (~AESL_inst_dft.temp_131_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_131_loc_channel_U.if_write) | (~AESL_inst_dft.temp_132_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_132_loc_channel_U.if_write) | (~AESL_inst_dft.temp_133_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_133_loc_channel_U.if_write) | (~AESL_inst_dft.temp_134_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_134_loc_channel_U.if_write) | (~AESL_inst_dft.temp_135_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_135_loc_channel_U.if_write) | (~AESL_inst_dft.temp_136_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_136_loc_channel_U.if_write) | (~AESL_inst_dft.temp_137_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_137_loc_channel_U.if_write) | (~AESL_inst_dft.temp_138_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_138_loc_channel_U.if_write) | (~AESL_inst_dft.temp_139_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_139_loc_channel_U.if_write) | (~AESL_inst_dft.temp_140_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_140_loc_channel_U.if_write) | (~AESL_inst_dft.temp_141_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_141_loc_channel_U.if_write) | (~AESL_inst_dft.temp_142_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_142_loc_channel_U.if_write) | (~AESL_inst_dft.temp_143_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_143_loc_channel_U.if_write) | (~AESL_inst_dft.temp_144_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_144_loc_channel_U.if_write) | (~AESL_inst_dft.temp_145_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_145_loc_channel_U.if_write) | (~AESL_inst_dft.temp_146_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_146_loc_channel_U.if_write) | (~AESL_inst_dft.temp_147_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_147_loc_channel_U.if_write) | (~AESL_inst_dft.temp_148_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_148_loc_channel_U.if_write) | (~AESL_inst_dft.temp_149_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_149_loc_channel_U.if_write) | (~AESL_inst_dft.temp_150_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_150_loc_channel_U.if_write) | (~AESL_inst_dft.temp_151_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_151_loc_channel_U.if_write) | (~AESL_inst_dft.temp_152_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_152_loc_channel_U.if_write) | (~AESL_inst_dft.temp_153_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_153_loc_channel_U.if_write) | (~AESL_inst_dft.temp_154_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_154_loc_channel_U.if_write) | (~AESL_inst_dft.temp_155_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_155_loc_channel_U.if_write) | (~AESL_inst_dft.temp_156_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_156_loc_channel_U.if_write) | (~AESL_inst_dft.temp_157_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_157_loc_channel_U.if_write) | (~AESL_inst_dft.temp_158_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_158_loc_channel_U.if_write) | (~AESL_inst_dft.temp_159_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_159_loc_channel_U.if_write) | (~AESL_inst_dft.temp_160_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_160_loc_channel_U.if_write) | (~AESL_inst_dft.temp_161_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_161_loc_channel_U.if_write) | (~AESL_inst_dft.temp_162_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_162_loc_channel_U.if_write) | (~AESL_inst_dft.temp_163_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_163_loc_channel_U.if_write) | (~AESL_inst_dft.temp_164_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_164_loc_channel_U.if_write) | (~AESL_inst_dft.temp_165_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_165_loc_channel_U.if_write) | (~AESL_inst_dft.temp_166_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_166_loc_channel_U.if_write) | (~AESL_inst_dft.temp_167_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_167_loc_channel_U.if_write) | (~AESL_inst_dft.temp_168_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_168_loc_channel_U.if_write) | (~AESL_inst_dft.temp_169_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_169_loc_channel_U.if_write) | (~AESL_inst_dft.temp_170_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_170_loc_channel_U.if_write) | (~AESL_inst_dft.temp_171_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_171_loc_channel_U.if_write) | (~AESL_inst_dft.temp_172_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_172_loc_channel_U.if_write) | (~AESL_inst_dft.temp_173_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_173_loc_channel_U.if_write) | (~AESL_inst_dft.temp_174_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_174_loc_channel_U.if_write) | (~AESL_inst_dft.temp_175_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_175_loc_channel_U.if_write) | (~AESL_inst_dft.temp_176_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_176_loc_channel_U.if_write) | (~AESL_inst_dft.temp_177_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_177_loc_channel_U.if_write) | (~AESL_inst_dft.temp_178_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_178_loc_channel_U.if_write) | (~AESL_inst_dft.temp_179_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_179_loc_channel_U.if_write) | (~AESL_inst_dft.temp_180_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_180_loc_channel_U.if_write) | (~AESL_inst_dft.temp_181_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_181_loc_channel_U.if_write) | (~AESL_inst_dft.temp_182_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_182_loc_channel_U.if_write) | (~AESL_inst_dft.temp_183_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_183_loc_channel_U.if_write) | (~AESL_inst_dft.temp_184_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_184_loc_channel_U.if_write) | (~AESL_inst_dft.temp_185_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_185_loc_channel_U.if_write) | (~AESL_inst_dft.temp_186_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_186_loc_channel_U.if_write) | (~AESL_inst_dft.temp_187_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_187_loc_channel_U.if_write) | (~AESL_inst_dft.temp_188_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_188_loc_channel_U.if_write) | (~AESL_inst_dft.temp_189_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_189_loc_channel_U.if_write) | (~AESL_inst_dft.temp_190_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_190_loc_channel_U.if_write) | (~AESL_inst_dft.temp_191_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_191_loc_channel_U.if_write) | (~AESL_inst_dft.temp_192_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_192_loc_channel_U.if_write) | (~AESL_inst_dft.temp_193_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_193_loc_channel_U.if_write) | (~AESL_inst_dft.temp_194_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_194_loc_channel_U.if_write) | (~AESL_inst_dft.temp_195_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_195_loc_channel_U.if_write) | (~AESL_inst_dft.temp_196_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_196_loc_channel_U.if_write) | (~AESL_inst_dft.temp_197_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_197_loc_channel_U.if_write) | (~AESL_inst_dft.temp_198_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_198_loc_channel_U.if_write) | (~AESL_inst_dft.temp_199_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_199_loc_channel_U.if_write) | (~AESL_inst_dft.temp_200_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_200_loc_channel_U.if_write) | (~AESL_inst_dft.temp_201_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_201_loc_channel_U.if_write) | (~AESL_inst_dft.temp_202_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_202_loc_channel_U.if_write) | (~AESL_inst_dft.temp_203_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_203_loc_channel_U.if_write) | (~AESL_inst_dft.temp_204_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_204_loc_channel_U.if_write) | (~AESL_inst_dft.temp_205_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_205_loc_channel_U.if_write) | (~AESL_inst_dft.temp_206_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_206_loc_channel_U.if_write) | (~AESL_inst_dft.temp_207_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_207_loc_channel_U.if_write) | (~AESL_inst_dft.temp_208_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_208_loc_channel_U.if_write) | (~AESL_inst_dft.temp_209_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_209_loc_channel_U.if_write) | (~AESL_inst_dft.temp_210_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_210_loc_channel_U.if_write) | (~AESL_inst_dft.temp_211_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_211_loc_channel_U.if_write) | (~AESL_inst_dft.temp_212_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_212_loc_channel_U.if_write) | (~AESL_inst_dft.temp_213_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_213_loc_channel_U.if_write) | (~AESL_inst_dft.temp_214_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_214_loc_channel_U.if_write) | (~AESL_inst_dft.temp_215_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_215_loc_channel_U.if_write) | (~AESL_inst_dft.temp_216_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_216_loc_channel_U.if_write) | (~AESL_inst_dft.temp_217_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_217_loc_channel_U.if_write) | (~AESL_inst_dft.temp_218_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_218_loc_channel_U.if_write) | (~AESL_inst_dft.temp_219_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_219_loc_channel_U.if_write) | (~AESL_inst_dft.temp_220_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_220_loc_channel_U.if_write) | (~AESL_inst_dft.temp_221_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_221_loc_channel_U.if_write) | (~AESL_inst_dft.temp_222_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_222_loc_channel_U.if_write) | (~AESL_inst_dft.temp_223_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_223_loc_channel_U.if_write) | (~AESL_inst_dft.temp_224_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_224_loc_channel_U.if_write) | (~AESL_inst_dft.temp_225_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_225_loc_channel_U.if_write) | (~AESL_inst_dft.temp_226_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_226_loc_channel_U.if_write) | (~AESL_inst_dft.temp_227_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_227_loc_channel_U.if_write) | (~AESL_inst_dft.temp_228_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_228_loc_channel_U.if_write) | (~AESL_inst_dft.temp_229_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_229_loc_channel_U.if_write) | (~AESL_inst_dft.temp_230_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_230_loc_channel_U.if_write) | (~AESL_inst_dft.temp_231_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_231_loc_channel_U.if_write) | (~AESL_inst_dft.temp_232_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_232_loc_channel_U.if_write) | (~AESL_inst_dft.temp_233_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_233_loc_channel_U.if_write) | (~AESL_inst_dft.temp_234_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_234_loc_channel_U.if_write) | (~AESL_inst_dft.temp_235_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_235_loc_channel_U.if_write) | (~AESL_inst_dft.temp_236_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_236_loc_channel_U.if_write) | (~AESL_inst_dft.temp_237_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_237_loc_channel_U.if_write) | (~AESL_inst_dft.temp_238_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_238_loc_channel_U.if_write) | (~AESL_inst_dft.temp_239_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_239_loc_channel_U.if_write) | (~AESL_inst_dft.temp_240_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_240_loc_channel_U.if_write) | (~AESL_inst_dft.temp_241_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_241_loc_channel_U.if_write) | (~AESL_inst_dft.temp_242_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_242_loc_channel_U.if_write) | (~AESL_inst_dft.temp_243_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_243_loc_channel_U.if_write) | (~AESL_inst_dft.temp_244_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_244_loc_channel_U.if_write) | (~AESL_inst_dft.temp_245_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_245_loc_channel_U.if_write) | (~AESL_inst_dft.temp_246_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_246_loc_channel_U.if_write) | (~AESL_inst_dft.temp_247_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_247_loc_channel_U.if_write) | (~AESL_inst_dft.temp_248_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_248_loc_channel_U.if_write) | (~AESL_inst_dft.temp_249_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_249_loc_channel_U.if_write) | (~AESL_inst_dft.temp_250_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_250_loc_channel_U.if_write) | (~AESL_inst_dft.temp_251_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_251_loc_channel_U.if_write) | (~AESL_inst_dft.temp_252_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_252_loc_channel_U.if_write) | (~AESL_inst_dft.temp_253_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_253_loc_channel_U.if_write) | (~AESL_inst_dft.temp_254_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_254_loc_channel_U.if_write) | (~AESL_inst_dft.temp_255_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_255_loc_channel_U.if_write);
    assign proc_1_input_sync_blk[0] = 1'b0 | (AESL_inst_dft.ap_sync_Loop_VITIS_LOOP_21_2_proc_U0_ap_ready & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.ap_sync_Loop_VITIS_LOOP_16_1_proc_U0_ap_ready);
    assign proc_1_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (proc_1_data_FIFO_blk[0] | proc_1_data_PIPO_blk[0] | proc_1_start_FIFO_blk[0] | proc_1_TLF_FIFO_blk[0] | proc_1_input_sync_blk[0] | proc_1_output_sync_blk[0]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[1 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[0];


    wire [1:0] dl_in_vec_comb = dl_in_vec & ~{1{all_finish}};
    AESL_deadlock_report_unit #(2) AESL_deadlock_report_unit_inst (
        .dl_reset(dl_reset),
        .dl_clock(dl_clock),
        .dl_in_vec(dl_in_vec_comb),
        .ap_done_reg_0(ap_done_reg_0),
        .dl_detect_out(dl_detect_out),
        .origin(origin),
        .token_clear(token_clear));

endmodule
