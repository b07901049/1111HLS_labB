`timescale 1 ns / 1 ps

module AESL_deadlock_report_unit #( parameter PROC_NUM = 4 ) (
    input dl_reset,
    input dl_clock,
    input [PROC_NUM - 1:0] dl_in_vec,
    input ap_done_reg_0,
    output dl_detect_out,
    output reg [PROC_NUM - 1:0] origin,
    output token_clear);
   
    // FSM states
    localparam ST_IDLE = 3'b000;
    localparam ST_FILTER_FAKE = 3'b001;
    localparam ST_DL_DETECTED = 3'b010;
    localparam ST_DL_REPORT = 3'b100;

    reg find_df_deadlock;
    reg [2:0] CS_fsm;
    reg [2:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    reg [31:0] dl_keep_cnt;
    integer i;
    integer fp;

    // FSM State machine
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end
    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg or dl_keep_cnt) begin
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_FILTER_FAKE;
                end
                else begin
                    NS_fsm = ST_IDLE;
                end
            end
            ST_FILTER_FAKE: begin
                if (dl_keep_cnt >= 32'd1000) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else if (dl_detect_reg != (dl_detect_reg & dl_in_vec)) begin
                    NS_fsm = ST_IDLE;
                end
                else begin
                    NS_fsm = ST_FILTER_FAKE;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if (dl_detect_reg != dl_done_reg) begin
                    NS_fsm = ST_DL_REPORT;
                end
                else begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            default: NS_fsm = ST_IDLE;
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_keep_cnt <= 32'h0;
        end
        else begin
            if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg == (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= dl_keep_cnt + 32'h1;
            end
            else if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg != (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= 32'h0;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = (|dl_detect_reg) && (CS_fsm == ST_DL_DETECTED || CS_fsm == ST_DL_REPORT);

    // dl_done_reg record the cycles has been reported
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    wire [PROC_NUM*PROC_NUM - 1:0] origin_tmp;
    assign origin_tmp[PROC_NUM - 1:0] = (dl_detect_reg[0] & ~dl_done_reg[0]) ? 'b1 : 'b0;
    genvar j;
    generate
    for(j = 1;j < PROC_NUM;j = j + 1) begin: F1
        assign origin_tmp[j*PROC_NUM +: PROC_NUM] = (dl_detect_reg[j] & ~dl_done_reg[j]) ? ('b1 << j) : origin_tmp[(j - 1)*PROC_NUM +: PROC_NUM];
    end
    endgenerate
    always @ (CS_fsm or origin_tmp) begin
        if (CS_fsm == ST_DL_DETECTED) begin
            origin = origin_tmp[(PROC_NUM - 1)*PROC_NUM +: PROC_NUM];
        end
        else begin
            origin = 'b0;
        end
    end

    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // find_df_deadlock to report the deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            find_df_deadlock <= 1'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED && dl_detect_reg == dl_done_reg) begin
                find_df_deadlock <= 1'b1;
            end
            else if (CS_fsm == ST_IDLE) begin
                find_df_deadlock <= 1'b0;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [336:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "dft.Loop_VITIS_LOOP_16_1_proc_U0";
                end
                1 : begin
                    proc_path = "dft.Loop_VITIS_LOOP_21_2_proc_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [336:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num, input integer record_time);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [336:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [288:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin
                    case(index2)
                    1: begin
                        if (AESL_inst_dft.ap_sync_Loop_VITIS_LOOP_16_1_proc_U0_ap_ready & AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_idle & ~AESL_inst_dft.ap_sync_Loop_VITIS_LOOP_21_2_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'dft.Loop_VITIS_LOOP_21_2_proc_U0'");
                        end
                    end
                    endcase
                end
                1 : begin
                    case(index2)
                    0: begin
                        if (~AESL_inst_dft.temp_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_1_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_1_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_1_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_1_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_1_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_1_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_1_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_1_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_2_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_2_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_2_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_2_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_2_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_2_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_2_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_2_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_3_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_3_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_3_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_3_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_3_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_3_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_3_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_3_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_4_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_4_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_4_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_4_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_4_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_4_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_4_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_4_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_5_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_5_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_5_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_5_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_5_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_5_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_5_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_5_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_6_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_6_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_6_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_6_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_6_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_6_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_6_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_6_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_7_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_7_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_7_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_7_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_7_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_7_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_7_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_7_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_8_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_8_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_8_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_8_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_8_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_8_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_8_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_8_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_9_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_9_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_9_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_9_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_9_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_9_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_9_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_9_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_10_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_10_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_10_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_10_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_10_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_10_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_10_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_10_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_11_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_11_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_11_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_11_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_11_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_11_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_11_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_11_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_12_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_12_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_12_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_12_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_12_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_12_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_12_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_12_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_13_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_13_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_13_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_13_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_13_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_13_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_13_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_13_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_14_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_14_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_14_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_14_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_14_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_14_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_14_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_14_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_15_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_15_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_15_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_15_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_15_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_15_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_15_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_15_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_16_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_16_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_16_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_16_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_16_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_16_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_16_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_16_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_17_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_17_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_17_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_17_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_17_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_17_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_17_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_17_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_18_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_18_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_18_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_18_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_18_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_18_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_18_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_18_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_19_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_19_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_19_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_19_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_19_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_19_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_19_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_19_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_20_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_20_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_20_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_20_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_20_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_20_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_20_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_20_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_21_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_21_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_21_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_21_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_21_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_21_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_21_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_21_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_22_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_22_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_22_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_22_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_22_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_22_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_22_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_22_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_23_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_23_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_23_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_23_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_23_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_23_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_23_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_23_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_24_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_24_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_24_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_24_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_24_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_24_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_24_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_24_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_25_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_25_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_25_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_25_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_25_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_25_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_25_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_25_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_26_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_26_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_26_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_26_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_26_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_26_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_26_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_26_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_27_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_27_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_27_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_27_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_27_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_27_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_27_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_27_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_28_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_28_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_28_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_28_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_28_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_28_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_28_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_28_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_29_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_29_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_29_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_29_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_29_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_29_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_29_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_29_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_30_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_30_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_30_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_30_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_30_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_30_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_30_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_30_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_31_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_31_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_31_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_31_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_31_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_31_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_31_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_31_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_32_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_32_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_32_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_32_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_32_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_32_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_32_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_32_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_33_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_33_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_33_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_33_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_33_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_33_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_33_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_33_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_34_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_34_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_34_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_34_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_34_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_34_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_34_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_34_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_35_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_35_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_35_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_35_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_35_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_35_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_35_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_35_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_36_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_36_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_36_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_36_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_36_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_36_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_36_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_36_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_37_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_37_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_37_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_37_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_37_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_37_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_37_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_37_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_38_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_38_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_38_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_38_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_38_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_38_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_38_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_38_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_39_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_39_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_39_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_39_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_39_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_39_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_39_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_39_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_40_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_40_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_40_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_40_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_40_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_40_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_40_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_40_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_41_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_41_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_41_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_41_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_41_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_41_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_41_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_41_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_42_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_42_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_42_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_42_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_42_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_42_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_42_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_42_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_43_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_43_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_43_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_43_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_43_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_43_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_43_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_43_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_44_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_44_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_44_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_44_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_44_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_44_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_44_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_44_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_45_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_45_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_45_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_45_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_45_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_45_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_45_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_45_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_46_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_46_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_46_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_46_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_46_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_46_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_46_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_46_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_47_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_47_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_47_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_47_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_47_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_47_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_47_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_47_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_48_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_48_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_48_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_48_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_48_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_48_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_48_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_48_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_49_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_49_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_49_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_49_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_49_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_49_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_49_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_49_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_50_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_50_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_50_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_50_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_50_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_50_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_50_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_50_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_51_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_51_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_51_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_51_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_51_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_51_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_51_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_51_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_52_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_52_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_52_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_52_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_52_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_52_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_52_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_52_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_53_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_53_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_53_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_53_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_53_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_53_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_53_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_53_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_54_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_54_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_54_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_54_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_54_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_54_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_54_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_54_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_55_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_55_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_55_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_55_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_55_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_55_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_55_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_55_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_56_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_56_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_56_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_56_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_56_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_56_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_56_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_56_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_57_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_57_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_57_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_57_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_57_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_57_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_57_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_57_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_58_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_58_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_58_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_58_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_58_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_58_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_58_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_58_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_59_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_59_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_59_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_59_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_59_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_59_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_59_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_59_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_60_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_60_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_60_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_60_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_60_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_60_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_60_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_60_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_61_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_61_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_61_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_61_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_61_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_61_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_61_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_61_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_62_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_62_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_62_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_62_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_62_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_62_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_62_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_62_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_63_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_63_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_63_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_63_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_63_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_63_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_63_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_63_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_64_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_64_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_64_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_64_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_64_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_64_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_64_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_64_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_65_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_65_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_65_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_65_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_65_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_65_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_65_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_65_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_66_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_66_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_66_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_66_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_66_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_66_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_66_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_66_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_67_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_67_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_67_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_67_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_67_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_67_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_67_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_67_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_68_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_68_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_68_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_68_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_68_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_68_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_68_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_68_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_69_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_69_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_69_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_69_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_69_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_69_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_69_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_69_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_70_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_70_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_70_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_70_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_70_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_70_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_70_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_70_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_71_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_71_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_71_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_71_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_71_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_71_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_71_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_71_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_72_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_72_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_72_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_72_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_72_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_72_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_72_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_72_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_73_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_73_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_73_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_73_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_73_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_73_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_73_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_73_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_74_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_74_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_74_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_74_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_74_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_74_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_74_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_74_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_75_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_75_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_75_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_75_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_75_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_75_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_75_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_75_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_76_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_76_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_76_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_76_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_76_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_76_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_76_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_76_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_77_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_77_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_77_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_77_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_77_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_77_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_77_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_77_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_78_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_78_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_78_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_78_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_78_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_78_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_78_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_78_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_79_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_79_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_79_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_79_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_79_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_79_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_79_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_79_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_80_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_80_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_80_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_80_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_80_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_80_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_80_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_80_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_81_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_81_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_81_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_81_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_81_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_81_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_81_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_81_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_82_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_82_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_82_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_82_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_82_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_82_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_82_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_82_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_83_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_83_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_83_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_83_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_83_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_83_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_83_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_83_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_84_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_84_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_84_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_84_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_84_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_84_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_84_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_84_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_85_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_85_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_85_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_85_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_85_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_85_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_85_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_85_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_86_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_86_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_86_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_86_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_86_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_86_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_86_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_86_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_87_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_87_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_87_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_87_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_87_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_87_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_87_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_87_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_88_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_88_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_88_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_88_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_88_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_88_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_88_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_88_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_89_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_89_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_89_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_89_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_89_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_89_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_89_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_89_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_90_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_90_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_90_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_90_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_90_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_90_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_90_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_90_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_91_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_91_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_91_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_91_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_91_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_91_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_91_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_91_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_92_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_92_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_92_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_92_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_92_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_92_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_92_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_92_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_93_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_93_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_93_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_93_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_93_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_93_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_93_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_93_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_94_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_94_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_94_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_94_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_94_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_94_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_94_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_94_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_95_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_95_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_95_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_95_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_95_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_95_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_95_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_95_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_96_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_96_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_96_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_96_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_96_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_96_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_96_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_96_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_97_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_97_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_97_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_97_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_97_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_97_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_97_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_97_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_98_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_98_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_98_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_98_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_98_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_98_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_98_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_98_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_99_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_99_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_99_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_99_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_99_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_99_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_99_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_99_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_100_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_100_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_100_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_100_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_100_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_100_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_100_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_100_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_101_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_101_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_101_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_101_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_101_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_101_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_101_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_101_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_102_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_102_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_102_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_102_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_102_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_102_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_102_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_102_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_103_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_103_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_103_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_103_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_103_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_103_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_103_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_103_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_104_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_104_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_104_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_104_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_104_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_104_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_104_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_104_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_105_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_105_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_105_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_105_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_105_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_105_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_105_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_105_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_106_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_106_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_106_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_106_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_106_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_106_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_106_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_106_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_107_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_107_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_107_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_107_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_107_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_107_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_107_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_107_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_108_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_108_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_108_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_108_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_108_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_108_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_108_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_108_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_109_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_109_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_109_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_109_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_109_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_109_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_109_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_109_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_110_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_110_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_110_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_110_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_110_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_110_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_110_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_110_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_111_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_111_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_111_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_111_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_111_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_111_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_111_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_111_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_112_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_112_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_112_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_112_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_112_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_112_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_112_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_112_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_113_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_113_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_113_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_113_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_113_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_113_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_113_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_113_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_114_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_114_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_114_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_114_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_114_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_114_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_114_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_114_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_115_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_115_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_115_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_115_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_115_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_115_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_115_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_115_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_116_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_116_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_116_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_116_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_116_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_116_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_116_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_116_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_117_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_117_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_117_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_117_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_117_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_117_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_117_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_117_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_118_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_118_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_118_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_118_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_118_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_118_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_118_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_118_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_119_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_119_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_119_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_119_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_119_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_119_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_119_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_119_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_120_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_120_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_120_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_120_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_120_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_120_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_120_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_120_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_121_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_121_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_121_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_121_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_121_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_121_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_121_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_121_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_122_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_122_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_122_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_122_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_122_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_122_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_122_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_122_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_123_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_123_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_123_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_123_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_123_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_123_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_123_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_123_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_124_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_124_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_124_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_124_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_124_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_124_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_124_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_124_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_125_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_125_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_125_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_125_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_125_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_125_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_125_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_125_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_126_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_126_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_126_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_126_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_126_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_126_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_126_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_126_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_127_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_127_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_127_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_127_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_127_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_127_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_127_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_127_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_128_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_128_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_128_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_128_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_128_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_128_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_128_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_128_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_129_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_129_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_129_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_129_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_129_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_129_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_129_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_129_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_130_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_130_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_130_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_130_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_130_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_130_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_130_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_130_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_131_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_131_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_131_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_131_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_131_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_131_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_131_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_131_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_132_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_132_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_132_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_132_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_132_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_132_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_132_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_132_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_133_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_133_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_133_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_133_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_133_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_133_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_133_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_133_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_134_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_134_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_134_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_134_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_134_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_134_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_134_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_134_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_135_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_135_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_135_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_135_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_135_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_135_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_135_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_135_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_136_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_136_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_136_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_136_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_136_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_136_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_136_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_136_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_137_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_137_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_137_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_137_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_137_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_137_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_137_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_137_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_138_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_138_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_138_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_138_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_138_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_138_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_138_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_138_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_139_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_139_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_139_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_139_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_139_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_139_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_139_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_139_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_140_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_140_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_140_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_140_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_140_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_140_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_140_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_140_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_141_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_141_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_141_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_141_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_141_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_141_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_141_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_141_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_142_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_142_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_142_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_142_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_142_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_142_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_142_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_142_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_143_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_143_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_143_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_143_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_143_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_143_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_143_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_143_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_144_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_144_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_144_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_144_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_144_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_144_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_144_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_144_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_145_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_145_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_145_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_145_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_145_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_145_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_145_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_145_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_146_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_146_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_146_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_146_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_146_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_146_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_146_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_146_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_147_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_147_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_147_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_147_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_147_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_147_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_147_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_147_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_148_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_148_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_148_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_148_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_148_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_148_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_148_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_148_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_149_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_149_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_149_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_149_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_149_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_149_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_149_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_149_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_150_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_150_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_150_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_150_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_150_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_150_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_150_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_150_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_151_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_151_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_151_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_151_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_151_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_151_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_151_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_151_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_152_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_152_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_152_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_152_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_152_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_152_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_152_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_152_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_153_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_153_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_153_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_153_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_153_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_153_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_153_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_153_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_154_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_154_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_154_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_154_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_154_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_154_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_154_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_154_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_155_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_155_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_155_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_155_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_155_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_155_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_155_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_155_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_156_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_156_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_156_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_156_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_156_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_156_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_156_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_156_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_157_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_157_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_157_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_157_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_157_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_157_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_157_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_157_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_158_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_158_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_158_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_158_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_158_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_158_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_158_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_158_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_159_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_159_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_159_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_159_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_159_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_159_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_159_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_159_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_160_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_160_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_160_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_160_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_160_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_160_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_160_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_160_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_161_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_161_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_161_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_161_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_161_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_161_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_161_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_161_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_162_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_162_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_162_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_162_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_162_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_162_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_162_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_162_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_163_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_163_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_163_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_163_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_163_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_163_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_163_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_163_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_164_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_164_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_164_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_164_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_164_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_164_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_164_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_164_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_165_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_165_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_165_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_165_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_165_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_165_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_165_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_165_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_166_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_166_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_166_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_166_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_166_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_166_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_166_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_166_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_167_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_167_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_167_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_167_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_167_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_167_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_167_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_167_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_168_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_168_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_168_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_168_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_168_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_168_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_168_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_168_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_169_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_169_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_169_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_169_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_169_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_169_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_169_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_169_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_170_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_170_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_170_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_170_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_170_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_170_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_170_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_170_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_171_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_171_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_171_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_171_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_171_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_171_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_171_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_171_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_172_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_172_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_172_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_172_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_172_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_172_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_172_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_172_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_173_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_173_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_173_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_173_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_173_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_173_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_173_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_173_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_174_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_174_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_174_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_174_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_174_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_174_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_174_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_174_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_175_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_175_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_175_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_175_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_175_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_175_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_175_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_175_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_176_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_176_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_176_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_176_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_176_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_176_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_176_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_176_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_177_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_177_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_177_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_177_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_177_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_177_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_177_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_177_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_178_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_178_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_178_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_178_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_178_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_178_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_178_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_178_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_179_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_179_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_179_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_179_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_179_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_179_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_179_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_179_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_180_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_180_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_180_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_180_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_180_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_180_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_180_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_180_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_181_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_181_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_181_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_181_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_181_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_181_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_181_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_181_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_182_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_182_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_182_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_182_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_182_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_182_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_182_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_182_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_183_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_183_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_183_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_183_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_183_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_183_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_183_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_183_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_184_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_184_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_184_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_184_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_184_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_184_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_184_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_184_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_185_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_185_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_185_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_185_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_185_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_185_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_185_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_185_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_186_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_186_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_186_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_186_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_186_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_186_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_186_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_186_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_187_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_187_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_187_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_187_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_187_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_187_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_187_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_187_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_188_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_188_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_188_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_188_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_188_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_188_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_188_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_188_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_189_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_189_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_189_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_189_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_189_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_189_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_189_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_189_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_190_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_190_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_190_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_190_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_190_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_190_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_190_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_190_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_191_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_191_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_191_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_191_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_191_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_191_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_191_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_191_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_192_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_192_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_192_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_192_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_192_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_192_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_192_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_192_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_193_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_193_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_193_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_193_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_193_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_193_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_193_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_193_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_194_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_194_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_194_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_194_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_194_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_194_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_194_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_194_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_195_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_195_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_195_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_195_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_195_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_195_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_195_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_195_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_196_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_196_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_196_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_196_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_196_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_196_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_196_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_196_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_197_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_197_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_197_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_197_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_197_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_197_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_197_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_197_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_198_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_198_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_198_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_198_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_198_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_198_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_198_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_198_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_199_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_199_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_199_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_199_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_199_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_199_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_199_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_199_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_200_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_200_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_200_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_200_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_200_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_200_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_200_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_200_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_201_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_201_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_201_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_201_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_201_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_201_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_201_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_201_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_202_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_202_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_202_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_202_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_202_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_202_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_202_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_202_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_203_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_203_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_203_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_203_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_203_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_203_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_203_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_203_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_204_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_204_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_204_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_204_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_204_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_204_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_204_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_204_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_205_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_205_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_205_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_205_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_205_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_205_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_205_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_205_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_206_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_206_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_206_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_206_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_206_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_206_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_206_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_206_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_207_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_207_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_207_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_207_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_207_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_207_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_207_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_207_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_208_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_208_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_208_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_208_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_208_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_208_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_208_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_208_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_209_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_209_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_209_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_209_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_209_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_209_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_209_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_209_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_210_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_210_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_210_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_210_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_210_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_210_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_210_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_210_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_211_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_211_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_211_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_211_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_211_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_211_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_211_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_211_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_212_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_212_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_212_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_212_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_212_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_212_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_212_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_212_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_213_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_213_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_213_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_213_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_213_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_213_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_213_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_213_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_214_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_214_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_214_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_214_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_214_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_214_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_214_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_214_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_215_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_215_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_215_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_215_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_215_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_215_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_215_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_215_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_216_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_216_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_216_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_216_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_216_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_216_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_216_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_216_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_217_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_217_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_217_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_217_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_217_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_217_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_217_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_217_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_218_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_218_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_218_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_218_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_218_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_218_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_218_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_218_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_219_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_219_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_219_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_219_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_219_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_219_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_219_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_219_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_220_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_220_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_220_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_220_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_220_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_220_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_220_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_220_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_221_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_221_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_221_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_221_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_221_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_221_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_221_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_221_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_222_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_222_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_222_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_222_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_222_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_222_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_222_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_222_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_223_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_223_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_223_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_223_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_223_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_223_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_223_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_223_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_224_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_224_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_224_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_224_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_224_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_224_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_224_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_224_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_225_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_225_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_225_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_225_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_225_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_225_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_225_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_225_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_226_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_226_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_226_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_226_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_226_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_226_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_226_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_226_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_227_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_227_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_227_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_227_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_227_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_227_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_227_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_227_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_228_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_228_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_228_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_228_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_228_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_228_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_228_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_228_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_229_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_229_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_229_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_229_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_229_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_229_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_229_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_229_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_230_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_230_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_230_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_230_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_230_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_230_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_230_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_230_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_231_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_231_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_231_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_231_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_231_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_231_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_231_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_231_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_232_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_232_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_232_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_232_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_232_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_232_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_232_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_232_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_233_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_233_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_233_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_233_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_233_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_233_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_233_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_233_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_234_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_234_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_234_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_234_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_234_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_234_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_234_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_234_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_235_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_235_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_235_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_235_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_235_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_235_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_235_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_235_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_236_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_236_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_236_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_236_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_236_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_236_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_236_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_236_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_237_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_237_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_237_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_237_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_237_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_237_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_237_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_237_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_238_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_238_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_238_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_238_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_238_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_238_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_238_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_238_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_239_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_239_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_239_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_239_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_239_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_239_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_239_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_239_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_240_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_240_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_240_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_240_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_240_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_240_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_240_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_240_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_241_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_241_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_241_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_241_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_241_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_241_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_241_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_241_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_242_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_242_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_242_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_242_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_242_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_242_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_242_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_242_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_243_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_243_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_243_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_243_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_243_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_243_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_243_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_243_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_244_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_244_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_244_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_244_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_244_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_244_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_244_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_244_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_245_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_245_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_245_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_245_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_245_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_245_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_245_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_245_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_246_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_246_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_246_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_246_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_246_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_246_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_246_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_246_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_247_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_247_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_247_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_247_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_247_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_247_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_247_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_247_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_248_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_248_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_248_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_248_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_248_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_248_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_248_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_248_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_249_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_249_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_249_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_249_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_249_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_249_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_249_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_249_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_250_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_250_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_250_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_250_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_250_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_250_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_250_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_250_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_251_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_251_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_251_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_251_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_251_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_251_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_251_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_251_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_252_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_252_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_252_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_252_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_252_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_252_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_252_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_252_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_253_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_253_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_253_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_253_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_253_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_253_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_253_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_253_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_254_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_254_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_254_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_254_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_254_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_254_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_254_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_254_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_dft.temp_255_loc_channel_U.if_empty_n & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.temp_255_loc_channel_U.if_write) begin
                            if (~AESL_inst_dft.temp_255_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'dft.temp_255_loc_channel_U' written by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_255_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_dft.temp_255_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'dft.temp_255_loc_channel_U' read by process 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path dft.temp_255_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (AESL_inst_dft.ap_sync_Loop_VITIS_LOOP_21_2_proc_U0_ap_ready & AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_idle & ~AESL_inst_dft.ap_sync_Loop_VITIS_LOOP_16_1_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'dft.Loop_VITIS_LOOP_16_1_proc_U0'");
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        integer record_time;
        wait (dl_reset == 1);
        cycle_id = 1;
        record_time = 0;
        while (1) begin
            @ (negedge dl_clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                            record_time = $time;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end((cycle_id - 1),record_time);
                        @(negedge dl_clock);
                        @(negedge dl_clock);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
endmodule
