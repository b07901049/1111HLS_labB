
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "df_fifo_interface.svh"
`include "df_fifo_monitor.svh"
`include "df_process_interface.svh"
`include "df_process_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);

    df_fifo_intf fifo_intf_1(clock,reset);
    assign fifo_intf_1.rd_en = AESL_inst_dft.temp_loc_channel_U.if_read & AESL_inst_dft.temp_loc_channel_U.if_empty_n;
    assign fifo_intf_1.wr_en = AESL_inst_dft.temp_loc_channel_U.if_write & AESL_inst_dft.temp_loc_channel_U.if_full_n;
    assign fifo_intf_1.fifo_rd_block = 0;
    assign fifo_intf_1.fifo_wr_block = 0;
    assign fifo_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_1;
    csv_file_dump cstatus_csv_dumper_1;
    df_fifo_monitor fifo_monitor_1;
    df_fifo_intf fifo_intf_2(clock,reset);
    assign fifo_intf_2.rd_en = AESL_inst_dft.temp_1_loc_channel_U.if_read & AESL_inst_dft.temp_1_loc_channel_U.if_empty_n;
    assign fifo_intf_2.wr_en = AESL_inst_dft.temp_1_loc_channel_U.if_write & AESL_inst_dft.temp_1_loc_channel_U.if_full_n;
    assign fifo_intf_2.fifo_rd_block = 0;
    assign fifo_intf_2.fifo_wr_block = 0;
    assign fifo_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_2;
    csv_file_dump cstatus_csv_dumper_2;
    df_fifo_monitor fifo_monitor_2;
    df_fifo_intf fifo_intf_3(clock,reset);
    assign fifo_intf_3.rd_en = AESL_inst_dft.temp_2_loc_channel_U.if_read & AESL_inst_dft.temp_2_loc_channel_U.if_empty_n;
    assign fifo_intf_3.wr_en = AESL_inst_dft.temp_2_loc_channel_U.if_write & AESL_inst_dft.temp_2_loc_channel_U.if_full_n;
    assign fifo_intf_3.fifo_rd_block = 0;
    assign fifo_intf_3.fifo_wr_block = 0;
    assign fifo_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_3;
    csv_file_dump cstatus_csv_dumper_3;
    df_fifo_monitor fifo_monitor_3;
    df_fifo_intf fifo_intf_4(clock,reset);
    assign fifo_intf_4.rd_en = AESL_inst_dft.temp_3_loc_channel_U.if_read & AESL_inst_dft.temp_3_loc_channel_U.if_empty_n;
    assign fifo_intf_4.wr_en = AESL_inst_dft.temp_3_loc_channel_U.if_write & AESL_inst_dft.temp_3_loc_channel_U.if_full_n;
    assign fifo_intf_4.fifo_rd_block = 0;
    assign fifo_intf_4.fifo_wr_block = 0;
    assign fifo_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_4;
    csv_file_dump cstatus_csv_dumper_4;
    df_fifo_monitor fifo_monitor_4;
    df_fifo_intf fifo_intf_5(clock,reset);
    assign fifo_intf_5.rd_en = AESL_inst_dft.temp_4_loc_channel_U.if_read & AESL_inst_dft.temp_4_loc_channel_U.if_empty_n;
    assign fifo_intf_5.wr_en = AESL_inst_dft.temp_4_loc_channel_U.if_write & AESL_inst_dft.temp_4_loc_channel_U.if_full_n;
    assign fifo_intf_5.fifo_rd_block = 0;
    assign fifo_intf_5.fifo_wr_block = 0;
    assign fifo_intf_5.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_5;
    csv_file_dump cstatus_csv_dumper_5;
    df_fifo_monitor fifo_monitor_5;
    df_fifo_intf fifo_intf_6(clock,reset);
    assign fifo_intf_6.rd_en = AESL_inst_dft.temp_5_loc_channel_U.if_read & AESL_inst_dft.temp_5_loc_channel_U.if_empty_n;
    assign fifo_intf_6.wr_en = AESL_inst_dft.temp_5_loc_channel_U.if_write & AESL_inst_dft.temp_5_loc_channel_U.if_full_n;
    assign fifo_intf_6.fifo_rd_block = 0;
    assign fifo_intf_6.fifo_wr_block = 0;
    assign fifo_intf_6.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_6;
    csv_file_dump cstatus_csv_dumper_6;
    df_fifo_monitor fifo_monitor_6;
    df_fifo_intf fifo_intf_7(clock,reset);
    assign fifo_intf_7.rd_en = AESL_inst_dft.temp_6_loc_channel_U.if_read & AESL_inst_dft.temp_6_loc_channel_U.if_empty_n;
    assign fifo_intf_7.wr_en = AESL_inst_dft.temp_6_loc_channel_U.if_write & AESL_inst_dft.temp_6_loc_channel_U.if_full_n;
    assign fifo_intf_7.fifo_rd_block = 0;
    assign fifo_intf_7.fifo_wr_block = 0;
    assign fifo_intf_7.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_7;
    csv_file_dump cstatus_csv_dumper_7;
    df_fifo_monitor fifo_monitor_7;
    df_fifo_intf fifo_intf_8(clock,reset);
    assign fifo_intf_8.rd_en = AESL_inst_dft.temp_7_loc_channel_U.if_read & AESL_inst_dft.temp_7_loc_channel_U.if_empty_n;
    assign fifo_intf_8.wr_en = AESL_inst_dft.temp_7_loc_channel_U.if_write & AESL_inst_dft.temp_7_loc_channel_U.if_full_n;
    assign fifo_intf_8.fifo_rd_block = 0;
    assign fifo_intf_8.fifo_wr_block = 0;
    assign fifo_intf_8.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_8;
    csv_file_dump cstatus_csv_dumper_8;
    df_fifo_monitor fifo_monitor_8;
    df_fifo_intf fifo_intf_9(clock,reset);
    assign fifo_intf_9.rd_en = AESL_inst_dft.temp_8_loc_channel_U.if_read & AESL_inst_dft.temp_8_loc_channel_U.if_empty_n;
    assign fifo_intf_9.wr_en = AESL_inst_dft.temp_8_loc_channel_U.if_write & AESL_inst_dft.temp_8_loc_channel_U.if_full_n;
    assign fifo_intf_9.fifo_rd_block = 0;
    assign fifo_intf_9.fifo_wr_block = 0;
    assign fifo_intf_9.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_9;
    csv_file_dump cstatus_csv_dumper_9;
    df_fifo_monitor fifo_monitor_9;
    df_fifo_intf fifo_intf_10(clock,reset);
    assign fifo_intf_10.rd_en = AESL_inst_dft.temp_9_loc_channel_U.if_read & AESL_inst_dft.temp_9_loc_channel_U.if_empty_n;
    assign fifo_intf_10.wr_en = AESL_inst_dft.temp_9_loc_channel_U.if_write & AESL_inst_dft.temp_9_loc_channel_U.if_full_n;
    assign fifo_intf_10.fifo_rd_block = 0;
    assign fifo_intf_10.fifo_wr_block = 0;
    assign fifo_intf_10.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_10;
    csv_file_dump cstatus_csv_dumper_10;
    df_fifo_monitor fifo_monitor_10;
    df_fifo_intf fifo_intf_11(clock,reset);
    assign fifo_intf_11.rd_en = AESL_inst_dft.temp_10_loc_channel_U.if_read & AESL_inst_dft.temp_10_loc_channel_U.if_empty_n;
    assign fifo_intf_11.wr_en = AESL_inst_dft.temp_10_loc_channel_U.if_write & AESL_inst_dft.temp_10_loc_channel_U.if_full_n;
    assign fifo_intf_11.fifo_rd_block = 0;
    assign fifo_intf_11.fifo_wr_block = 0;
    assign fifo_intf_11.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_11;
    csv_file_dump cstatus_csv_dumper_11;
    df_fifo_monitor fifo_monitor_11;
    df_fifo_intf fifo_intf_12(clock,reset);
    assign fifo_intf_12.rd_en = AESL_inst_dft.temp_11_loc_channel_U.if_read & AESL_inst_dft.temp_11_loc_channel_U.if_empty_n;
    assign fifo_intf_12.wr_en = AESL_inst_dft.temp_11_loc_channel_U.if_write & AESL_inst_dft.temp_11_loc_channel_U.if_full_n;
    assign fifo_intf_12.fifo_rd_block = 0;
    assign fifo_intf_12.fifo_wr_block = 0;
    assign fifo_intf_12.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_12;
    csv_file_dump cstatus_csv_dumper_12;
    df_fifo_monitor fifo_monitor_12;
    df_fifo_intf fifo_intf_13(clock,reset);
    assign fifo_intf_13.rd_en = AESL_inst_dft.temp_12_loc_channel_U.if_read & AESL_inst_dft.temp_12_loc_channel_U.if_empty_n;
    assign fifo_intf_13.wr_en = AESL_inst_dft.temp_12_loc_channel_U.if_write & AESL_inst_dft.temp_12_loc_channel_U.if_full_n;
    assign fifo_intf_13.fifo_rd_block = 0;
    assign fifo_intf_13.fifo_wr_block = 0;
    assign fifo_intf_13.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_13;
    csv_file_dump cstatus_csv_dumper_13;
    df_fifo_monitor fifo_monitor_13;
    df_fifo_intf fifo_intf_14(clock,reset);
    assign fifo_intf_14.rd_en = AESL_inst_dft.temp_13_loc_channel_U.if_read & AESL_inst_dft.temp_13_loc_channel_U.if_empty_n;
    assign fifo_intf_14.wr_en = AESL_inst_dft.temp_13_loc_channel_U.if_write & AESL_inst_dft.temp_13_loc_channel_U.if_full_n;
    assign fifo_intf_14.fifo_rd_block = 0;
    assign fifo_intf_14.fifo_wr_block = 0;
    assign fifo_intf_14.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_14;
    csv_file_dump cstatus_csv_dumper_14;
    df_fifo_monitor fifo_monitor_14;
    df_fifo_intf fifo_intf_15(clock,reset);
    assign fifo_intf_15.rd_en = AESL_inst_dft.temp_14_loc_channel_U.if_read & AESL_inst_dft.temp_14_loc_channel_U.if_empty_n;
    assign fifo_intf_15.wr_en = AESL_inst_dft.temp_14_loc_channel_U.if_write & AESL_inst_dft.temp_14_loc_channel_U.if_full_n;
    assign fifo_intf_15.fifo_rd_block = 0;
    assign fifo_intf_15.fifo_wr_block = 0;
    assign fifo_intf_15.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_15;
    csv_file_dump cstatus_csv_dumper_15;
    df_fifo_monitor fifo_monitor_15;
    df_fifo_intf fifo_intf_16(clock,reset);
    assign fifo_intf_16.rd_en = AESL_inst_dft.temp_15_loc_channel_U.if_read & AESL_inst_dft.temp_15_loc_channel_U.if_empty_n;
    assign fifo_intf_16.wr_en = AESL_inst_dft.temp_15_loc_channel_U.if_write & AESL_inst_dft.temp_15_loc_channel_U.if_full_n;
    assign fifo_intf_16.fifo_rd_block = 0;
    assign fifo_intf_16.fifo_wr_block = 0;
    assign fifo_intf_16.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_16;
    csv_file_dump cstatus_csv_dumper_16;
    df_fifo_monitor fifo_monitor_16;
    df_fifo_intf fifo_intf_17(clock,reset);
    assign fifo_intf_17.rd_en = AESL_inst_dft.temp_16_loc_channel_U.if_read & AESL_inst_dft.temp_16_loc_channel_U.if_empty_n;
    assign fifo_intf_17.wr_en = AESL_inst_dft.temp_16_loc_channel_U.if_write & AESL_inst_dft.temp_16_loc_channel_U.if_full_n;
    assign fifo_intf_17.fifo_rd_block = 0;
    assign fifo_intf_17.fifo_wr_block = 0;
    assign fifo_intf_17.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_17;
    csv_file_dump cstatus_csv_dumper_17;
    df_fifo_monitor fifo_monitor_17;
    df_fifo_intf fifo_intf_18(clock,reset);
    assign fifo_intf_18.rd_en = AESL_inst_dft.temp_17_loc_channel_U.if_read & AESL_inst_dft.temp_17_loc_channel_U.if_empty_n;
    assign fifo_intf_18.wr_en = AESL_inst_dft.temp_17_loc_channel_U.if_write & AESL_inst_dft.temp_17_loc_channel_U.if_full_n;
    assign fifo_intf_18.fifo_rd_block = 0;
    assign fifo_intf_18.fifo_wr_block = 0;
    assign fifo_intf_18.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_18;
    csv_file_dump cstatus_csv_dumper_18;
    df_fifo_monitor fifo_monitor_18;
    df_fifo_intf fifo_intf_19(clock,reset);
    assign fifo_intf_19.rd_en = AESL_inst_dft.temp_18_loc_channel_U.if_read & AESL_inst_dft.temp_18_loc_channel_U.if_empty_n;
    assign fifo_intf_19.wr_en = AESL_inst_dft.temp_18_loc_channel_U.if_write & AESL_inst_dft.temp_18_loc_channel_U.if_full_n;
    assign fifo_intf_19.fifo_rd_block = 0;
    assign fifo_intf_19.fifo_wr_block = 0;
    assign fifo_intf_19.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_19;
    csv_file_dump cstatus_csv_dumper_19;
    df_fifo_monitor fifo_monitor_19;
    df_fifo_intf fifo_intf_20(clock,reset);
    assign fifo_intf_20.rd_en = AESL_inst_dft.temp_19_loc_channel_U.if_read & AESL_inst_dft.temp_19_loc_channel_U.if_empty_n;
    assign fifo_intf_20.wr_en = AESL_inst_dft.temp_19_loc_channel_U.if_write & AESL_inst_dft.temp_19_loc_channel_U.if_full_n;
    assign fifo_intf_20.fifo_rd_block = 0;
    assign fifo_intf_20.fifo_wr_block = 0;
    assign fifo_intf_20.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_20;
    csv_file_dump cstatus_csv_dumper_20;
    df_fifo_monitor fifo_monitor_20;
    df_fifo_intf fifo_intf_21(clock,reset);
    assign fifo_intf_21.rd_en = AESL_inst_dft.temp_20_loc_channel_U.if_read & AESL_inst_dft.temp_20_loc_channel_U.if_empty_n;
    assign fifo_intf_21.wr_en = AESL_inst_dft.temp_20_loc_channel_U.if_write & AESL_inst_dft.temp_20_loc_channel_U.if_full_n;
    assign fifo_intf_21.fifo_rd_block = 0;
    assign fifo_intf_21.fifo_wr_block = 0;
    assign fifo_intf_21.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_21;
    csv_file_dump cstatus_csv_dumper_21;
    df_fifo_monitor fifo_monitor_21;
    df_fifo_intf fifo_intf_22(clock,reset);
    assign fifo_intf_22.rd_en = AESL_inst_dft.temp_21_loc_channel_U.if_read & AESL_inst_dft.temp_21_loc_channel_U.if_empty_n;
    assign fifo_intf_22.wr_en = AESL_inst_dft.temp_21_loc_channel_U.if_write & AESL_inst_dft.temp_21_loc_channel_U.if_full_n;
    assign fifo_intf_22.fifo_rd_block = 0;
    assign fifo_intf_22.fifo_wr_block = 0;
    assign fifo_intf_22.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_22;
    csv_file_dump cstatus_csv_dumper_22;
    df_fifo_monitor fifo_monitor_22;
    df_fifo_intf fifo_intf_23(clock,reset);
    assign fifo_intf_23.rd_en = AESL_inst_dft.temp_22_loc_channel_U.if_read & AESL_inst_dft.temp_22_loc_channel_U.if_empty_n;
    assign fifo_intf_23.wr_en = AESL_inst_dft.temp_22_loc_channel_U.if_write & AESL_inst_dft.temp_22_loc_channel_U.if_full_n;
    assign fifo_intf_23.fifo_rd_block = 0;
    assign fifo_intf_23.fifo_wr_block = 0;
    assign fifo_intf_23.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_23;
    csv_file_dump cstatus_csv_dumper_23;
    df_fifo_monitor fifo_monitor_23;
    df_fifo_intf fifo_intf_24(clock,reset);
    assign fifo_intf_24.rd_en = AESL_inst_dft.temp_23_loc_channel_U.if_read & AESL_inst_dft.temp_23_loc_channel_U.if_empty_n;
    assign fifo_intf_24.wr_en = AESL_inst_dft.temp_23_loc_channel_U.if_write & AESL_inst_dft.temp_23_loc_channel_U.if_full_n;
    assign fifo_intf_24.fifo_rd_block = 0;
    assign fifo_intf_24.fifo_wr_block = 0;
    assign fifo_intf_24.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_24;
    csv_file_dump cstatus_csv_dumper_24;
    df_fifo_monitor fifo_monitor_24;
    df_fifo_intf fifo_intf_25(clock,reset);
    assign fifo_intf_25.rd_en = AESL_inst_dft.temp_24_loc_channel_U.if_read & AESL_inst_dft.temp_24_loc_channel_U.if_empty_n;
    assign fifo_intf_25.wr_en = AESL_inst_dft.temp_24_loc_channel_U.if_write & AESL_inst_dft.temp_24_loc_channel_U.if_full_n;
    assign fifo_intf_25.fifo_rd_block = 0;
    assign fifo_intf_25.fifo_wr_block = 0;
    assign fifo_intf_25.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_25;
    csv_file_dump cstatus_csv_dumper_25;
    df_fifo_monitor fifo_monitor_25;
    df_fifo_intf fifo_intf_26(clock,reset);
    assign fifo_intf_26.rd_en = AESL_inst_dft.temp_25_loc_channel_U.if_read & AESL_inst_dft.temp_25_loc_channel_U.if_empty_n;
    assign fifo_intf_26.wr_en = AESL_inst_dft.temp_25_loc_channel_U.if_write & AESL_inst_dft.temp_25_loc_channel_U.if_full_n;
    assign fifo_intf_26.fifo_rd_block = 0;
    assign fifo_intf_26.fifo_wr_block = 0;
    assign fifo_intf_26.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_26;
    csv_file_dump cstatus_csv_dumper_26;
    df_fifo_monitor fifo_monitor_26;
    df_fifo_intf fifo_intf_27(clock,reset);
    assign fifo_intf_27.rd_en = AESL_inst_dft.temp_26_loc_channel_U.if_read & AESL_inst_dft.temp_26_loc_channel_U.if_empty_n;
    assign fifo_intf_27.wr_en = AESL_inst_dft.temp_26_loc_channel_U.if_write & AESL_inst_dft.temp_26_loc_channel_U.if_full_n;
    assign fifo_intf_27.fifo_rd_block = 0;
    assign fifo_intf_27.fifo_wr_block = 0;
    assign fifo_intf_27.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_27;
    csv_file_dump cstatus_csv_dumper_27;
    df_fifo_monitor fifo_monitor_27;
    df_fifo_intf fifo_intf_28(clock,reset);
    assign fifo_intf_28.rd_en = AESL_inst_dft.temp_27_loc_channel_U.if_read & AESL_inst_dft.temp_27_loc_channel_U.if_empty_n;
    assign fifo_intf_28.wr_en = AESL_inst_dft.temp_27_loc_channel_U.if_write & AESL_inst_dft.temp_27_loc_channel_U.if_full_n;
    assign fifo_intf_28.fifo_rd_block = 0;
    assign fifo_intf_28.fifo_wr_block = 0;
    assign fifo_intf_28.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_28;
    csv_file_dump cstatus_csv_dumper_28;
    df_fifo_monitor fifo_monitor_28;
    df_fifo_intf fifo_intf_29(clock,reset);
    assign fifo_intf_29.rd_en = AESL_inst_dft.temp_28_loc_channel_U.if_read & AESL_inst_dft.temp_28_loc_channel_U.if_empty_n;
    assign fifo_intf_29.wr_en = AESL_inst_dft.temp_28_loc_channel_U.if_write & AESL_inst_dft.temp_28_loc_channel_U.if_full_n;
    assign fifo_intf_29.fifo_rd_block = 0;
    assign fifo_intf_29.fifo_wr_block = 0;
    assign fifo_intf_29.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_29;
    csv_file_dump cstatus_csv_dumper_29;
    df_fifo_monitor fifo_monitor_29;
    df_fifo_intf fifo_intf_30(clock,reset);
    assign fifo_intf_30.rd_en = AESL_inst_dft.temp_29_loc_channel_U.if_read & AESL_inst_dft.temp_29_loc_channel_U.if_empty_n;
    assign fifo_intf_30.wr_en = AESL_inst_dft.temp_29_loc_channel_U.if_write & AESL_inst_dft.temp_29_loc_channel_U.if_full_n;
    assign fifo_intf_30.fifo_rd_block = 0;
    assign fifo_intf_30.fifo_wr_block = 0;
    assign fifo_intf_30.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_30;
    csv_file_dump cstatus_csv_dumper_30;
    df_fifo_monitor fifo_monitor_30;
    df_fifo_intf fifo_intf_31(clock,reset);
    assign fifo_intf_31.rd_en = AESL_inst_dft.temp_30_loc_channel_U.if_read & AESL_inst_dft.temp_30_loc_channel_U.if_empty_n;
    assign fifo_intf_31.wr_en = AESL_inst_dft.temp_30_loc_channel_U.if_write & AESL_inst_dft.temp_30_loc_channel_U.if_full_n;
    assign fifo_intf_31.fifo_rd_block = 0;
    assign fifo_intf_31.fifo_wr_block = 0;
    assign fifo_intf_31.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_31;
    csv_file_dump cstatus_csv_dumper_31;
    df_fifo_monitor fifo_monitor_31;
    df_fifo_intf fifo_intf_32(clock,reset);
    assign fifo_intf_32.rd_en = AESL_inst_dft.temp_31_loc_channel_U.if_read & AESL_inst_dft.temp_31_loc_channel_U.if_empty_n;
    assign fifo_intf_32.wr_en = AESL_inst_dft.temp_31_loc_channel_U.if_write & AESL_inst_dft.temp_31_loc_channel_U.if_full_n;
    assign fifo_intf_32.fifo_rd_block = 0;
    assign fifo_intf_32.fifo_wr_block = 0;
    assign fifo_intf_32.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_32;
    csv_file_dump cstatus_csv_dumper_32;
    df_fifo_monitor fifo_monitor_32;
    df_fifo_intf fifo_intf_33(clock,reset);
    assign fifo_intf_33.rd_en = AESL_inst_dft.temp_32_loc_channel_U.if_read & AESL_inst_dft.temp_32_loc_channel_U.if_empty_n;
    assign fifo_intf_33.wr_en = AESL_inst_dft.temp_32_loc_channel_U.if_write & AESL_inst_dft.temp_32_loc_channel_U.if_full_n;
    assign fifo_intf_33.fifo_rd_block = 0;
    assign fifo_intf_33.fifo_wr_block = 0;
    assign fifo_intf_33.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_33;
    csv_file_dump cstatus_csv_dumper_33;
    df_fifo_monitor fifo_monitor_33;
    df_fifo_intf fifo_intf_34(clock,reset);
    assign fifo_intf_34.rd_en = AESL_inst_dft.temp_33_loc_channel_U.if_read & AESL_inst_dft.temp_33_loc_channel_U.if_empty_n;
    assign fifo_intf_34.wr_en = AESL_inst_dft.temp_33_loc_channel_U.if_write & AESL_inst_dft.temp_33_loc_channel_U.if_full_n;
    assign fifo_intf_34.fifo_rd_block = 0;
    assign fifo_intf_34.fifo_wr_block = 0;
    assign fifo_intf_34.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_34;
    csv_file_dump cstatus_csv_dumper_34;
    df_fifo_monitor fifo_monitor_34;
    df_fifo_intf fifo_intf_35(clock,reset);
    assign fifo_intf_35.rd_en = AESL_inst_dft.temp_34_loc_channel_U.if_read & AESL_inst_dft.temp_34_loc_channel_U.if_empty_n;
    assign fifo_intf_35.wr_en = AESL_inst_dft.temp_34_loc_channel_U.if_write & AESL_inst_dft.temp_34_loc_channel_U.if_full_n;
    assign fifo_intf_35.fifo_rd_block = 0;
    assign fifo_intf_35.fifo_wr_block = 0;
    assign fifo_intf_35.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_35;
    csv_file_dump cstatus_csv_dumper_35;
    df_fifo_monitor fifo_monitor_35;
    df_fifo_intf fifo_intf_36(clock,reset);
    assign fifo_intf_36.rd_en = AESL_inst_dft.temp_35_loc_channel_U.if_read & AESL_inst_dft.temp_35_loc_channel_U.if_empty_n;
    assign fifo_intf_36.wr_en = AESL_inst_dft.temp_35_loc_channel_U.if_write & AESL_inst_dft.temp_35_loc_channel_U.if_full_n;
    assign fifo_intf_36.fifo_rd_block = 0;
    assign fifo_intf_36.fifo_wr_block = 0;
    assign fifo_intf_36.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_36;
    csv_file_dump cstatus_csv_dumper_36;
    df_fifo_monitor fifo_monitor_36;
    df_fifo_intf fifo_intf_37(clock,reset);
    assign fifo_intf_37.rd_en = AESL_inst_dft.temp_36_loc_channel_U.if_read & AESL_inst_dft.temp_36_loc_channel_U.if_empty_n;
    assign fifo_intf_37.wr_en = AESL_inst_dft.temp_36_loc_channel_U.if_write & AESL_inst_dft.temp_36_loc_channel_U.if_full_n;
    assign fifo_intf_37.fifo_rd_block = 0;
    assign fifo_intf_37.fifo_wr_block = 0;
    assign fifo_intf_37.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_37;
    csv_file_dump cstatus_csv_dumper_37;
    df_fifo_monitor fifo_monitor_37;
    df_fifo_intf fifo_intf_38(clock,reset);
    assign fifo_intf_38.rd_en = AESL_inst_dft.temp_37_loc_channel_U.if_read & AESL_inst_dft.temp_37_loc_channel_U.if_empty_n;
    assign fifo_intf_38.wr_en = AESL_inst_dft.temp_37_loc_channel_U.if_write & AESL_inst_dft.temp_37_loc_channel_U.if_full_n;
    assign fifo_intf_38.fifo_rd_block = 0;
    assign fifo_intf_38.fifo_wr_block = 0;
    assign fifo_intf_38.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_38;
    csv_file_dump cstatus_csv_dumper_38;
    df_fifo_monitor fifo_monitor_38;
    df_fifo_intf fifo_intf_39(clock,reset);
    assign fifo_intf_39.rd_en = AESL_inst_dft.temp_38_loc_channel_U.if_read & AESL_inst_dft.temp_38_loc_channel_U.if_empty_n;
    assign fifo_intf_39.wr_en = AESL_inst_dft.temp_38_loc_channel_U.if_write & AESL_inst_dft.temp_38_loc_channel_U.if_full_n;
    assign fifo_intf_39.fifo_rd_block = 0;
    assign fifo_intf_39.fifo_wr_block = 0;
    assign fifo_intf_39.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_39;
    csv_file_dump cstatus_csv_dumper_39;
    df_fifo_monitor fifo_monitor_39;
    df_fifo_intf fifo_intf_40(clock,reset);
    assign fifo_intf_40.rd_en = AESL_inst_dft.temp_39_loc_channel_U.if_read & AESL_inst_dft.temp_39_loc_channel_U.if_empty_n;
    assign fifo_intf_40.wr_en = AESL_inst_dft.temp_39_loc_channel_U.if_write & AESL_inst_dft.temp_39_loc_channel_U.if_full_n;
    assign fifo_intf_40.fifo_rd_block = 0;
    assign fifo_intf_40.fifo_wr_block = 0;
    assign fifo_intf_40.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_40;
    csv_file_dump cstatus_csv_dumper_40;
    df_fifo_monitor fifo_monitor_40;
    df_fifo_intf fifo_intf_41(clock,reset);
    assign fifo_intf_41.rd_en = AESL_inst_dft.temp_40_loc_channel_U.if_read & AESL_inst_dft.temp_40_loc_channel_U.if_empty_n;
    assign fifo_intf_41.wr_en = AESL_inst_dft.temp_40_loc_channel_U.if_write & AESL_inst_dft.temp_40_loc_channel_U.if_full_n;
    assign fifo_intf_41.fifo_rd_block = 0;
    assign fifo_intf_41.fifo_wr_block = 0;
    assign fifo_intf_41.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_41;
    csv_file_dump cstatus_csv_dumper_41;
    df_fifo_monitor fifo_monitor_41;
    df_fifo_intf fifo_intf_42(clock,reset);
    assign fifo_intf_42.rd_en = AESL_inst_dft.temp_41_loc_channel_U.if_read & AESL_inst_dft.temp_41_loc_channel_U.if_empty_n;
    assign fifo_intf_42.wr_en = AESL_inst_dft.temp_41_loc_channel_U.if_write & AESL_inst_dft.temp_41_loc_channel_U.if_full_n;
    assign fifo_intf_42.fifo_rd_block = 0;
    assign fifo_intf_42.fifo_wr_block = 0;
    assign fifo_intf_42.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_42;
    csv_file_dump cstatus_csv_dumper_42;
    df_fifo_monitor fifo_monitor_42;
    df_fifo_intf fifo_intf_43(clock,reset);
    assign fifo_intf_43.rd_en = AESL_inst_dft.temp_42_loc_channel_U.if_read & AESL_inst_dft.temp_42_loc_channel_U.if_empty_n;
    assign fifo_intf_43.wr_en = AESL_inst_dft.temp_42_loc_channel_U.if_write & AESL_inst_dft.temp_42_loc_channel_U.if_full_n;
    assign fifo_intf_43.fifo_rd_block = 0;
    assign fifo_intf_43.fifo_wr_block = 0;
    assign fifo_intf_43.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_43;
    csv_file_dump cstatus_csv_dumper_43;
    df_fifo_monitor fifo_monitor_43;
    df_fifo_intf fifo_intf_44(clock,reset);
    assign fifo_intf_44.rd_en = AESL_inst_dft.temp_43_loc_channel_U.if_read & AESL_inst_dft.temp_43_loc_channel_U.if_empty_n;
    assign fifo_intf_44.wr_en = AESL_inst_dft.temp_43_loc_channel_U.if_write & AESL_inst_dft.temp_43_loc_channel_U.if_full_n;
    assign fifo_intf_44.fifo_rd_block = 0;
    assign fifo_intf_44.fifo_wr_block = 0;
    assign fifo_intf_44.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_44;
    csv_file_dump cstatus_csv_dumper_44;
    df_fifo_monitor fifo_monitor_44;
    df_fifo_intf fifo_intf_45(clock,reset);
    assign fifo_intf_45.rd_en = AESL_inst_dft.temp_44_loc_channel_U.if_read & AESL_inst_dft.temp_44_loc_channel_U.if_empty_n;
    assign fifo_intf_45.wr_en = AESL_inst_dft.temp_44_loc_channel_U.if_write & AESL_inst_dft.temp_44_loc_channel_U.if_full_n;
    assign fifo_intf_45.fifo_rd_block = 0;
    assign fifo_intf_45.fifo_wr_block = 0;
    assign fifo_intf_45.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_45;
    csv_file_dump cstatus_csv_dumper_45;
    df_fifo_monitor fifo_monitor_45;
    df_fifo_intf fifo_intf_46(clock,reset);
    assign fifo_intf_46.rd_en = AESL_inst_dft.temp_45_loc_channel_U.if_read & AESL_inst_dft.temp_45_loc_channel_U.if_empty_n;
    assign fifo_intf_46.wr_en = AESL_inst_dft.temp_45_loc_channel_U.if_write & AESL_inst_dft.temp_45_loc_channel_U.if_full_n;
    assign fifo_intf_46.fifo_rd_block = 0;
    assign fifo_intf_46.fifo_wr_block = 0;
    assign fifo_intf_46.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_46;
    csv_file_dump cstatus_csv_dumper_46;
    df_fifo_monitor fifo_monitor_46;
    df_fifo_intf fifo_intf_47(clock,reset);
    assign fifo_intf_47.rd_en = AESL_inst_dft.temp_46_loc_channel_U.if_read & AESL_inst_dft.temp_46_loc_channel_U.if_empty_n;
    assign fifo_intf_47.wr_en = AESL_inst_dft.temp_46_loc_channel_U.if_write & AESL_inst_dft.temp_46_loc_channel_U.if_full_n;
    assign fifo_intf_47.fifo_rd_block = 0;
    assign fifo_intf_47.fifo_wr_block = 0;
    assign fifo_intf_47.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_47;
    csv_file_dump cstatus_csv_dumper_47;
    df_fifo_monitor fifo_monitor_47;
    df_fifo_intf fifo_intf_48(clock,reset);
    assign fifo_intf_48.rd_en = AESL_inst_dft.temp_47_loc_channel_U.if_read & AESL_inst_dft.temp_47_loc_channel_U.if_empty_n;
    assign fifo_intf_48.wr_en = AESL_inst_dft.temp_47_loc_channel_U.if_write & AESL_inst_dft.temp_47_loc_channel_U.if_full_n;
    assign fifo_intf_48.fifo_rd_block = 0;
    assign fifo_intf_48.fifo_wr_block = 0;
    assign fifo_intf_48.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_48;
    csv_file_dump cstatus_csv_dumper_48;
    df_fifo_monitor fifo_monitor_48;
    df_fifo_intf fifo_intf_49(clock,reset);
    assign fifo_intf_49.rd_en = AESL_inst_dft.temp_48_loc_channel_U.if_read & AESL_inst_dft.temp_48_loc_channel_U.if_empty_n;
    assign fifo_intf_49.wr_en = AESL_inst_dft.temp_48_loc_channel_U.if_write & AESL_inst_dft.temp_48_loc_channel_U.if_full_n;
    assign fifo_intf_49.fifo_rd_block = 0;
    assign fifo_intf_49.fifo_wr_block = 0;
    assign fifo_intf_49.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_49;
    csv_file_dump cstatus_csv_dumper_49;
    df_fifo_monitor fifo_monitor_49;
    df_fifo_intf fifo_intf_50(clock,reset);
    assign fifo_intf_50.rd_en = AESL_inst_dft.temp_49_loc_channel_U.if_read & AESL_inst_dft.temp_49_loc_channel_U.if_empty_n;
    assign fifo_intf_50.wr_en = AESL_inst_dft.temp_49_loc_channel_U.if_write & AESL_inst_dft.temp_49_loc_channel_U.if_full_n;
    assign fifo_intf_50.fifo_rd_block = 0;
    assign fifo_intf_50.fifo_wr_block = 0;
    assign fifo_intf_50.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_50;
    csv_file_dump cstatus_csv_dumper_50;
    df_fifo_monitor fifo_monitor_50;
    df_fifo_intf fifo_intf_51(clock,reset);
    assign fifo_intf_51.rd_en = AESL_inst_dft.temp_50_loc_channel_U.if_read & AESL_inst_dft.temp_50_loc_channel_U.if_empty_n;
    assign fifo_intf_51.wr_en = AESL_inst_dft.temp_50_loc_channel_U.if_write & AESL_inst_dft.temp_50_loc_channel_U.if_full_n;
    assign fifo_intf_51.fifo_rd_block = 0;
    assign fifo_intf_51.fifo_wr_block = 0;
    assign fifo_intf_51.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_51;
    csv_file_dump cstatus_csv_dumper_51;
    df_fifo_monitor fifo_monitor_51;
    df_fifo_intf fifo_intf_52(clock,reset);
    assign fifo_intf_52.rd_en = AESL_inst_dft.temp_51_loc_channel_U.if_read & AESL_inst_dft.temp_51_loc_channel_U.if_empty_n;
    assign fifo_intf_52.wr_en = AESL_inst_dft.temp_51_loc_channel_U.if_write & AESL_inst_dft.temp_51_loc_channel_U.if_full_n;
    assign fifo_intf_52.fifo_rd_block = 0;
    assign fifo_intf_52.fifo_wr_block = 0;
    assign fifo_intf_52.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_52;
    csv_file_dump cstatus_csv_dumper_52;
    df_fifo_monitor fifo_monitor_52;
    df_fifo_intf fifo_intf_53(clock,reset);
    assign fifo_intf_53.rd_en = AESL_inst_dft.temp_52_loc_channel_U.if_read & AESL_inst_dft.temp_52_loc_channel_U.if_empty_n;
    assign fifo_intf_53.wr_en = AESL_inst_dft.temp_52_loc_channel_U.if_write & AESL_inst_dft.temp_52_loc_channel_U.if_full_n;
    assign fifo_intf_53.fifo_rd_block = 0;
    assign fifo_intf_53.fifo_wr_block = 0;
    assign fifo_intf_53.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_53;
    csv_file_dump cstatus_csv_dumper_53;
    df_fifo_monitor fifo_monitor_53;
    df_fifo_intf fifo_intf_54(clock,reset);
    assign fifo_intf_54.rd_en = AESL_inst_dft.temp_53_loc_channel_U.if_read & AESL_inst_dft.temp_53_loc_channel_U.if_empty_n;
    assign fifo_intf_54.wr_en = AESL_inst_dft.temp_53_loc_channel_U.if_write & AESL_inst_dft.temp_53_loc_channel_U.if_full_n;
    assign fifo_intf_54.fifo_rd_block = 0;
    assign fifo_intf_54.fifo_wr_block = 0;
    assign fifo_intf_54.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_54;
    csv_file_dump cstatus_csv_dumper_54;
    df_fifo_monitor fifo_monitor_54;
    df_fifo_intf fifo_intf_55(clock,reset);
    assign fifo_intf_55.rd_en = AESL_inst_dft.temp_54_loc_channel_U.if_read & AESL_inst_dft.temp_54_loc_channel_U.if_empty_n;
    assign fifo_intf_55.wr_en = AESL_inst_dft.temp_54_loc_channel_U.if_write & AESL_inst_dft.temp_54_loc_channel_U.if_full_n;
    assign fifo_intf_55.fifo_rd_block = 0;
    assign fifo_intf_55.fifo_wr_block = 0;
    assign fifo_intf_55.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_55;
    csv_file_dump cstatus_csv_dumper_55;
    df_fifo_monitor fifo_monitor_55;
    df_fifo_intf fifo_intf_56(clock,reset);
    assign fifo_intf_56.rd_en = AESL_inst_dft.temp_55_loc_channel_U.if_read & AESL_inst_dft.temp_55_loc_channel_U.if_empty_n;
    assign fifo_intf_56.wr_en = AESL_inst_dft.temp_55_loc_channel_U.if_write & AESL_inst_dft.temp_55_loc_channel_U.if_full_n;
    assign fifo_intf_56.fifo_rd_block = 0;
    assign fifo_intf_56.fifo_wr_block = 0;
    assign fifo_intf_56.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_56;
    csv_file_dump cstatus_csv_dumper_56;
    df_fifo_monitor fifo_monitor_56;
    df_fifo_intf fifo_intf_57(clock,reset);
    assign fifo_intf_57.rd_en = AESL_inst_dft.temp_56_loc_channel_U.if_read & AESL_inst_dft.temp_56_loc_channel_U.if_empty_n;
    assign fifo_intf_57.wr_en = AESL_inst_dft.temp_56_loc_channel_U.if_write & AESL_inst_dft.temp_56_loc_channel_U.if_full_n;
    assign fifo_intf_57.fifo_rd_block = 0;
    assign fifo_intf_57.fifo_wr_block = 0;
    assign fifo_intf_57.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_57;
    csv_file_dump cstatus_csv_dumper_57;
    df_fifo_monitor fifo_monitor_57;
    df_fifo_intf fifo_intf_58(clock,reset);
    assign fifo_intf_58.rd_en = AESL_inst_dft.temp_57_loc_channel_U.if_read & AESL_inst_dft.temp_57_loc_channel_U.if_empty_n;
    assign fifo_intf_58.wr_en = AESL_inst_dft.temp_57_loc_channel_U.if_write & AESL_inst_dft.temp_57_loc_channel_U.if_full_n;
    assign fifo_intf_58.fifo_rd_block = 0;
    assign fifo_intf_58.fifo_wr_block = 0;
    assign fifo_intf_58.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_58;
    csv_file_dump cstatus_csv_dumper_58;
    df_fifo_monitor fifo_monitor_58;
    df_fifo_intf fifo_intf_59(clock,reset);
    assign fifo_intf_59.rd_en = AESL_inst_dft.temp_58_loc_channel_U.if_read & AESL_inst_dft.temp_58_loc_channel_U.if_empty_n;
    assign fifo_intf_59.wr_en = AESL_inst_dft.temp_58_loc_channel_U.if_write & AESL_inst_dft.temp_58_loc_channel_U.if_full_n;
    assign fifo_intf_59.fifo_rd_block = 0;
    assign fifo_intf_59.fifo_wr_block = 0;
    assign fifo_intf_59.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_59;
    csv_file_dump cstatus_csv_dumper_59;
    df_fifo_monitor fifo_monitor_59;
    df_fifo_intf fifo_intf_60(clock,reset);
    assign fifo_intf_60.rd_en = AESL_inst_dft.temp_59_loc_channel_U.if_read & AESL_inst_dft.temp_59_loc_channel_U.if_empty_n;
    assign fifo_intf_60.wr_en = AESL_inst_dft.temp_59_loc_channel_U.if_write & AESL_inst_dft.temp_59_loc_channel_U.if_full_n;
    assign fifo_intf_60.fifo_rd_block = 0;
    assign fifo_intf_60.fifo_wr_block = 0;
    assign fifo_intf_60.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_60;
    csv_file_dump cstatus_csv_dumper_60;
    df_fifo_monitor fifo_monitor_60;
    df_fifo_intf fifo_intf_61(clock,reset);
    assign fifo_intf_61.rd_en = AESL_inst_dft.temp_60_loc_channel_U.if_read & AESL_inst_dft.temp_60_loc_channel_U.if_empty_n;
    assign fifo_intf_61.wr_en = AESL_inst_dft.temp_60_loc_channel_U.if_write & AESL_inst_dft.temp_60_loc_channel_U.if_full_n;
    assign fifo_intf_61.fifo_rd_block = 0;
    assign fifo_intf_61.fifo_wr_block = 0;
    assign fifo_intf_61.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_61;
    csv_file_dump cstatus_csv_dumper_61;
    df_fifo_monitor fifo_monitor_61;
    df_fifo_intf fifo_intf_62(clock,reset);
    assign fifo_intf_62.rd_en = AESL_inst_dft.temp_61_loc_channel_U.if_read & AESL_inst_dft.temp_61_loc_channel_U.if_empty_n;
    assign fifo_intf_62.wr_en = AESL_inst_dft.temp_61_loc_channel_U.if_write & AESL_inst_dft.temp_61_loc_channel_U.if_full_n;
    assign fifo_intf_62.fifo_rd_block = 0;
    assign fifo_intf_62.fifo_wr_block = 0;
    assign fifo_intf_62.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_62;
    csv_file_dump cstatus_csv_dumper_62;
    df_fifo_monitor fifo_monitor_62;
    df_fifo_intf fifo_intf_63(clock,reset);
    assign fifo_intf_63.rd_en = AESL_inst_dft.temp_62_loc_channel_U.if_read & AESL_inst_dft.temp_62_loc_channel_U.if_empty_n;
    assign fifo_intf_63.wr_en = AESL_inst_dft.temp_62_loc_channel_U.if_write & AESL_inst_dft.temp_62_loc_channel_U.if_full_n;
    assign fifo_intf_63.fifo_rd_block = 0;
    assign fifo_intf_63.fifo_wr_block = 0;
    assign fifo_intf_63.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_63;
    csv_file_dump cstatus_csv_dumper_63;
    df_fifo_monitor fifo_monitor_63;
    df_fifo_intf fifo_intf_64(clock,reset);
    assign fifo_intf_64.rd_en = AESL_inst_dft.temp_63_loc_channel_U.if_read & AESL_inst_dft.temp_63_loc_channel_U.if_empty_n;
    assign fifo_intf_64.wr_en = AESL_inst_dft.temp_63_loc_channel_U.if_write & AESL_inst_dft.temp_63_loc_channel_U.if_full_n;
    assign fifo_intf_64.fifo_rd_block = 0;
    assign fifo_intf_64.fifo_wr_block = 0;
    assign fifo_intf_64.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_64;
    csv_file_dump cstatus_csv_dumper_64;
    df_fifo_monitor fifo_monitor_64;
    df_fifo_intf fifo_intf_65(clock,reset);
    assign fifo_intf_65.rd_en = AESL_inst_dft.temp_64_loc_channel_U.if_read & AESL_inst_dft.temp_64_loc_channel_U.if_empty_n;
    assign fifo_intf_65.wr_en = AESL_inst_dft.temp_64_loc_channel_U.if_write & AESL_inst_dft.temp_64_loc_channel_U.if_full_n;
    assign fifo_intf_65.fifo_rd_block = 0;
    assign fifo_intf_65.fifo_wr_block = 0;
    assign fifo_intf_65.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_65;
    csv_file_dump cstatus_csv_dumper_65;
    df_fifo_monitor fifo_monitor_65;
    df_fifo_intf fifo_intf_66(clock,reset);
    assign fifo_intf_66.rd_en = AESL_inst_dft.temp_65_loc_channel_U.if_read & AESL_inst_dft.temp_65_loc_channel_U.if_empty_n;
    assign fifo_intf_66.wr_en = AESL_inst_dft.temp_65_loc_channel_U.if_write & AESL_inst_dft.temp_65_loc_channel_U.if_full_n;
    assign fifo_intf_66.fifo_rd_block = 0;
    assign fifo_intf_66.fifo_wr_block = 0;
    assign fifo_intf_66.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_66;
    csv_file_dump cstatus_csv_dumper_66;
    df_fifo_monitor fifo_monitor_66;
    df_fifo_intf fifo_intf_67(clock,reset);
    assign fifo_intf_67.rd_en = AESL_inst_dft.temp_66_loc_channel_U.if_read & AESL_inst_dft.temp_66_loc_channel_U.if_empty_n;
    assign fifo_intf_67.wr_en = AESL_inst_dft.temp_66_loc_channel_U.if_write & AESL_inst_dft.temp_66_loc_channel_U.if_full_n;
    assign fifo_intf_67.fifo_rd_block = 0;
    assign fifo_intf_67.fifo_wr_block = 0;
    assign fifo_intf_67.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_67;
    csv_file_dump cstatus_csv_dumper_67;
    df_fifo_monitor fifo_monitor_67;
    df_fifo_intf fifo_intf_68(clock,reset);
    assign fifo_intf_68.rd_en = AESL_inst_dft.temp_67_loc_channel_U.if_read & AESL_inst_dft.temp_67_loc_channel_U.if_empty_n;
    assign fifo_intf_68.wr_en = AESL_inst_dft.temp_67_loc_channel_U.if_write & AESL_inst_dft.temp_67_loc_channel_U.if_full_n;
    assign fifo_intf_68.fifo_rd_block = 0;
    assign fifo_intf_68.fifo_wr_block = 0;
    assign fifo_intf_68.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_68;
    csv_file_dump cstatus_csv_dumper_68;
    df_fifo_monitor fifo_monitor_68;
    df_fifo_intf fifo_intf_69(clock,reset);
    assign fifo_intf_69.rd_en = AESL_inst_dft.temp_68_loc_channel_U.if_read & AESL_inst_dft.temp_68_loc_channel_U.if_empty_n;
    assign fifo_intf_69.wr_en = AESL_inst_dft.temp_68_loc_channel_U.if_write & AESL_inst_dft.temp_68_loc_channel_U.if_full_n;
    assign fifo_intf_69.fifo_rd_block = 0;
    assign fifo_intf_69.fifo_wr_block = 0;
    assign fifo_intf_69.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_69;
    csv_file_dump cstatus_csv_dumper_69;
    df_fifo_monitor fifo_monitor_69;
    df_fifo_intf fifo_intf_70(clock,reset);
    assign fifo_intf_70.rd_en = AESL_inst_dft.temp_69_loc_channel_U.if_read & AESL_inst_dft.temp_69_loc_channel_U.if_empty_n;
    assign fifo_intf_70.wr_en = AESL_inst_dft.temp_69_loc_channel_U.if_write & AESL_inst_dft.temp_69_loc_channel_U.if_full_n;
    assign fifo_intf_70.fifo_rd_block = 0;
    assign fifo_intf_70.fifo_wr_block = 0;
    assign fifo_intf_70.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_70;
    csv_file_dump cstatus_csv_dumper_70;
    df_fifo_monitor fifo_monitor_70;
    df_fifo_intf fifo_intf_71(clock,reset);
    assign fifo_intf_71.rd_en = AESL_inst_dft.temp_70_loc_channel_U.if_read & AESL_inst_dft.temp_70_loc_channel_U.if_empty_n;
    assign fifo_intf_71.wr_en = AESL_inst_dft.temp_70_loc_channel_U.if_write & AESL_inst_dft.temp_70_loc_channel_U.if_full_n;
    assign fifo_intf_71.fifo_rd_block = 0;
    assign fifo_intf_71.fifo_wr_block = 0;
    assign fifo_intf_71.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_71;
    csv_file_dump cstatus_csv_dumper_71;
    df_fifo_monitor fifo_monitor_71;
    df_fifo_intf fifo_intf_72(clock,reset);
    assign fifo_intf_72.rd_en = AESL_inst_dft.temp_71_loc_channel_U.if_read & AESL_inst_dft.temp_71_loc_channel_U.if_empty_n;
    assign fifo_intf_72.wr_en = AESL_inst_dft.temp_71_loc_channel_U.if_write & AESL_inst_dft.temp_71_loc_channel_U.if_full_n;
    assign fifo_intf_72.fifo_rd_block = 0;
    assign fifo_intf_72.fifo_wr_block = 0;
    assign fifo_intf_72.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_72;
    csv_file_dump cstatus_csv_dumper_72;
    df_fifo_monitor fifo_monitor_72;
    df_fifo_intf fifo_intf_73(clock,reset);
    assign fifo_intf_73.rd_en = AESL_inst_dft.temp_72_loc_channel_U.if_read & AESL_inst_dft.temp_72_loc_channel_U.if_empty_n;
    assign fifo_intf_73.wr_en = AESL_inst_dft.temp_72_loc_channel_U.if_write & AESL_inst_dft.temp_72_loc_channel_U.if_full_n;
    assign fifo_intf_73.fifo_rd_block = 0;
    assign fifo_intf_73.fifo_wr_block = 0;
    assign fifo_intf_73.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_73;
    csv_file_dump cstatus_csv_dumper_73;
    df_fifo_monitor fifo_monitor_73;
    df_fifo_intf fifo_intf_74(clock,reset);
    assign fifo_intf_74.rd_en = AESL_inst_dft.temp_73_loc_channel_U.if_read & AESL_inst_dft.temp_73_loc_channel_U.if_empty_n;
    assign fifo_intf_74.wr_en = AESL_inst_dft.temp_73_loc_channel_U.if_write & AESL_inst_dft.temp_73_loc_channel_U.if_full_n;
    assign fifo_intf_74.fifo_rd_block = 0;
    assign fifo_intf_74.fifo_wr_block = 0;
    assign fifo_intf_74.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_74;
    csv_file_dump cstatus_csv_dumper_74;
    df_fifo_monitor fifo_monitor_74;
    df_fifo_intf fifo_intf_75(clock,reset);
    assign fifo_intf_75.rd_en = AESL_inst_dft.temp_74_loc_channel_U.if_read & AESL_inst_dft.temp_74_loc_channel_U.if_empty_n;
    assign fifo_intf_75.wr_en = AESL_inst_dft.temp_74_loc_channel_U.if_write & AESL_inst_dft.temp_74_loc_channel_U.if_full_n;
    assign fifo_intf_75.fifo_rd_block = 0;
    assign fifo_intf_75.fifo_wr_block = 0;
    assign fifo_intf_75.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_75;
    csv_file_dump cstatus_csv_dumper_75;
    df_fifo_monitor fifo_monitor_75;
    df_fifo_intf fifo_intf_76(clock,reset);
    assign fifo_intf_76.rd_en = AESL_inst_dft.temp_75_loc_channel_U.if_read & AESL_inst_dft.temp_75_loc_channel_U.if_empty_n;
    assign fifo_intf_76.wr_en = AESL_inst_dft.temp_75_loc_channel_U.if_write & AESL_inst_dft.temp_75_loc_channel_U.if_full_n;
    assign fifo_intf_76.fifo_rd_block = 0;
    assign fifo_intf_76.fifo_wr_block = 0;
    assign fifo_intf_76.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_76;
    csv_file_dump cstatus_csv_dumper_76;
    df_fifo_monitor fifo_monitor_76;
    df_fifo_intf fifo_intf_77(clock,reset);
    assign fifo_intf_77.rd_en = AESL_inst_dft.temp_76_loc_channel_U.if_read & AESL_inst_dft.temp_76_loc_channel_U.if_empty_n;
    assign fifo_intf_77.wr_en = AESL_inst_dft.temp_76_loc_channel_U.if_write & AESL_inst_dft.temp_76_loc_channel_U.if_full_n;
    assign fifo_intf_77.fifo_rd_block = 0;
    assign fifo_intf_77.fifo_wr_block = 0;
    assign fifo_intf_77.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_77;
    csv_file_dump cstatus_csv_dumper_77;
    df_fifo_monitor fifo_monitor_77;
    df_fifo_intf fifo_intf_78(clock,reset);
    assign fifo_intf_78.rd_en = AESL_inst_dft.temp_77_loc_channel_U.if_read & AESL_inst_dft.temp_77_loc_channel_U.if_empty_n;
    assign fifo_intf_78.wr_en = AESL_inst_dft.temp_77_loc_channel_U.if_write & AESL_inst_dft.temp_77_loc_channel_U.if_full_n;
    assign fifo_intf_78.fifo_rd_block = 0;
    assign fifo_intf_78.fifo_wr_block = 0;
    assign fifo_intf_78.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_78;
    csv_file_dump cstatus_csv_dumper_78;
    df_fifo_monitor fifo_monitor_78;
    df_fifo_intf fifo_intf_79(clock,reset);
    assign fifo_intf_79.rd_en = AESL_inst_dft.temp_78_loc_channel_U.if_read & AESL_inst_dft.temp_78_loc_channel_U.if_empty_n;
    assign fifo_intf_79.wr_en = AESL_inst_dft.temp_78_loc_channel_U.if_write & AESL_inst_dft.temp_78_loc_channel_U.if_full_n;
    assign fifo_intf_79.fifo_rd_block = 0;
    assign fifo_intf_79.fifo_wr_block = 0;
    assign fifo_intf_79.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_79;
    csv_file_dump cstatus_csv_dumper_79;
    df_fifo_monitor fifo_monitor_79;
    df_fifo_intf fifo_intf_80(clock,reset);
    assign fifo_intf_80.rd_en = AESL_inst_dft.temp_79_loc_channel_U.if_read & AESL_inst_dft.temp_79_loc_channel_U.if_empty_n;
    assign fifo_intf_80.wr_en = AESL_inst_dft.temp_79_loc_channel_U.if_write & AESL_inst_dft.temp_79_loc_channel_U.if_full_n;
    assign fifo_intf_80.fifo_rd_block = 0;
    assign fifo_intf_80.fifo_wr_block = 0;
    assign fifo_intf_80.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_80;
    csv_file_dump cstatus_csv_dumper_80;
    df_fifo_monitor fifo_monitor_80;
    df_fifo_intf fifo_intf_81(clock,reset);
    assign fifo_intf_81.rd_en = AESL_inst_dft.temp_80_loc_channel_U.if_read & AESL_inst_dft.temp_80_loc_channel_U.if_empty_n;
    assign fifo_intf_81.wr_en = AESL_inst_dft.temp_80_loc_channel_U.if_write & AESL_inst_dft.temp_80_loc_channel_U.if_full_n;
    assign fifo_intf_81.fifo_rd_block = 0;
    assign fifo_intf_81.fifo_wr_block = 0;
    assign fifo_intf_81.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_81;
    csv_file_dump cstatus_csv_dumper_81;
    df_fifo_monitor fifo_monitor_81;
    df_fifo_intf fifo_intf_82(clock,reset);
    assign fifo_intf_82.rd_en = AESL_inst_dft.temp_81_loc_channel_U.if_read & AESL_inst_dft.temp_81_loc_channel_U.if_empty_n;
    assign fifo_intf_82.wr_en = AESL_inst_dft.temp_81_loc_channel_U.if_write & AESL_inst_dft.temp_81_loc_channel_U.if_full_n;
    assign fifo_intf_82.fifo_rd_block = 0;
    assign fifo_intf_82.fifo_wr_block = 0;
    assign fifo_intf_82.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_82;
    csv_file_dump cstatus_csv_dumper_82;
    df_fifo_monitor fifo_monitor_82;
    df_fifo_intf fifo_intf_83(clock,reset);
    assign fifo_intf_83.rd_en = AESL_inst_dft.temp_82_loc_channel_U.if_read & AESL_inst_dft.temp_82_loc_channel_U.if_empty_n;
    assign fifo_intf_83.wr_en = AESL_inst_dft.temp_82_loc_channel_U.if_write & AESL_inst_dft.temp_82_loc_channel_U.if_full_n;
    assign fifo_intf_83.fifo_rd_block = 0;
    assign fifo_intf_83.fifo_wr_block = 0;
    assign fifo_intf_83.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_83;
    csv_file_dump cstatus_csv_dumper_83;
    df_fifo_monitor fifo_monitor_83;
    df_fifo_intf fifo_intf_84(clock,reset);
    assign fifo_intf_84.rd_en = AESL_inst_dft.temp_83_loc_channel_U.if_read & AESL_inst_dft.temp_83_loc_channel_U.if_empty_n;
    assign fifo_intf_84.wr_en = AESL_inst_dft.temp_83_loc_channel_U.if_write & AESL_inst_dft.temp_83_loc_channel_U.if_full_n;
    assign fifo_intf_84.fifo_rd_block = 0;
    assign fifo_intf_84.fifo_wr_block = 0;
    assign fifo_intf_84.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_84;
    csv_file_dump cstatus_csv_dumper_84;
    df_fifo_monitor fifo_monitor_84;
    df_fifo_intf fifo_intf_85(clock,reset);
    assign fifo_intf_85.rd_en = AESL_inst_dft.temp_84_loc_channel_U.if_read & AESL_inst_dft.temp_84_loc_channel_U.if_empty_n;
    assign fifo_intf_85.wr_en = AESL_inst_dft.temp_84_loc_channel_U.if_write & AESL_inst_dft.temp_84_loc_channel_U.if_full_n;
    assign fifo_intf_85.fifo_rd_block = 0;
    assign fifo_intf_85.fifo_wr_block = 0;
    assign fifo_intf_85.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_85;
    csv_file_dump cstatus_csv_dumper_85;
    df_fifo_monitor fifo_monitor_85;
    df_fifo_intf fifo_intf_86(clock,reset);
    assign fifo_intf_86.rd_en = AESL_inst_dft.temp_85_loc_channel_U.if_read & AESL_inst_dft.temp_85_loc_channel_U.if_empty_n;
    assign fifo_intf_86.wr_en = AESL_inst_dft.temp_85_loc_channel_U.if_write & AESL_inst_dft.temp_85_loc_channel_U.if_full_n;
    assign fifo_intf_86.fifo_rd_block = 0;
    assign fifo_intf_86.fifo_wr_block = 0;
    assign fifo_intf_86.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_86;
    csv_file_dump cstatus_csv_dumper_86;
    df_fifo_monitor fifo_monitor_86;
    df_fifo_intf fifo_intf_87(clock,reset);
    assign fifo_intf_87.rd_en = AESL_inst_dft.temp_86_loc_channel_U.if_read & AESL_inst_dft.temp_86_loc_channel_U.if_empty_n;
    assign fifo_intf_87.wr_en = AESL_inst_dft.temp_86_loc_channel_U.if_write & AESL_inst_dft.temp_86_loc_channel_U.if_full_n;
    assign fifo_intf_87.fifo_rd_block = 0;
    assign fifo_intf_87.fifo_wr_block = 0;
    assign fifo_intf_87.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_87;
    csv_file_dump cstatus_csv_dumper_87;
    df_fifo_monitor fifo_monitor_87;
    df_fifo_intf fifo_intf_88(clock,reset);
    assign fifo_intf_88.rd_en = AESL_inst_dft.temp_87_loc_channel_U.if_read & AESL_inst_dft.temp_87_loc_channel_U.if_empty_n;
    assign fifo_intf_88.wr_en = AESL_inst_dft.temp_87_loc_channel_U.if_write & AESL_inst_dft.temp_87_loc_channel_U.if_full_n;
    assign fifo_intf_88.fifo_rd_block = 0;
    assign fifo_intf_88.fifo_wr_block = 0;
    assign fifo_intf_88.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_88;
    csv_file_dump cstatus_csv_dumper_88;
    df_fifo_monitor fifo_monitor_88;
    df_fifo_intf fifo_intf_89(clock,reset);
    assign fifo_intf_89.rd_en = AESL_inst_dft.temp_88_loc_channel_U.if_read & AESL_inst_dft.temp_88_loc_channel_U.if_empty_n;
    assign fifo_intf_89.wr_en = AESL_inst_dft.temp_88_loc_channel_U.if_write & AESL_inst_dft.temp_88_loc_channel_U.if_full_n;
    assign fifo_intf_89.fifo_rd_block = 0;
    assign fifo_intf_89.fifo_wr_block = 0;
    assign fifo_intf_89.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_89;
    csv_file_dump cstatus_csv_dumper_89;
    df_fifo_monitor fifo_monitor_89;
    df_fifo_intf fifo_intf_90(clock,reset);
    assign fifo_intf_90.rd_en = AESL_inst_dft.temp_89_loc_channel_U.if_read & AESL_inst_dft.temp_89_loc_channel_U.if_empty_n;
    assign fifo_intf_90.wr_en = AESL_inst_dft.temp_89_loc_channel_U.if_write & AESL_inst_dft.temp_89_loc_channel_U.if_full_n;
    assign fifo_intf_90.fifo_rd_block = 0;
    assign fifo_intf_90.fifo_wr_block = 0;
    assign fifo_intf_90.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_90;
    csv_file_dump cstatus_csv_dumper_90;
    df_fifo_monitor fifo_monitor_90;
    df_fifo_intf fifo_intf_91(clock,reset);
    assign fifo_intf_91.rd_en = AESL_inst_dft.temp_90_loc_channel_U.if_read & AESL_inst_dft.temp_90_loc_channel_U.if_empty_n;
    assign fifo_intf_91.wr_en = AESL_inst_dft.temp_90_loc_channel_U.if_write & AESL_inst_dft.temp_90_loc_channel_U.if_full_n;
    assign fifo_intf_91.fifo_rd_block = 0;
    assign fifo_intf_91.fifo_wr_block = 0;
    assign fifo_intf_91.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_91;
    csv_file_dump cstatus_csv_dumper_91;
    df_fifo_monitor fifo_monitor_91;
    df_fifo_intf fifo_intf_92(clock,reset);
    assign fifo_intf_92.rd_en = AESL_inst_dft.temp_91_loc_channel_U.if_read & AESL_inst_dft.temp_91_loc_channel_U.if_empty_n;
    assign fifo_intf_92.wr_en = AESL_inst_dft.temp_91_loc_channel_U.if_write & AESL_inst_dft.temp_91_loc_channel_U.if_full_n;
    assign fifo_intf_92.fifo_rd_block = 0;
    assign fifo_intf_92.fifo_wr_block = 0;
    assign fifo_intf_92.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_92;
    csv_file_dump cstatus_csv_dumper_92;
    df_fifo_monitor fifo_monitor_92;
    df_fifo_intf fifo_intf_93(clock,reset);
    assign fifo_intf_93.rd_en = AESL_inst_dft.temp_92_loc_channel_U.if_read & AESL_inst_dft.temp_92_loc_channel_U.if_empty_n;
    assign fifo_intf_93.wr_en = AESL_inst_dft.temp_92_loc_channel_U.if_write & AESL_inst_dft.temp_92_loc_channel_U.if_full_n;
    assign fifo_intf_93.fifo_rd_block = 0;
    assign fifo_intf_93.fifo_wr_block = 0;
    assign fifo_intf_93.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_93;
    csv_file_dump cstatus_csv_dumper_93;
    df_fifo_monitor fifo_monitor_93;
    df_fifo_intf fifo_intf_94(clock,reset);
    assign fifo_intf_94.rd_en = AESL_inst_dft.temp_93_loc_channel_U.if_read & AESL_inst_dft.temp_93_loc_channel_U.if_empty_n;
    assign fifo_intf_94.wr_en = AESL_inst_dft.temp_93_loc_channel_U.if_write & AESL_inst_dft.temp_93_loc_channel_U.if_full_n;
    assign fifo_intf_94.fifo_rd_block = 0;
    assign fifo_intf_94.fifo_wr_block = 0;
    assign fifo_intf_94.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_94;
    csv_file_dump cstatus_csv_dumper_94;
    df_fifo_monitor fifo_monitor_94;
    df_fifo_intf fifo_intf_95(clock,reset);
    assign fifo_intf_95.rd_en = AESL_inst_dft.temp_94_loc_channel_U.if_read & AESL_inst_dft.temp_94_loc_channel_U.if_empty_n;
    assign fifo_intf_95.wr_en = AESL_inst_dft.temp_94_loc_channel_U.if_write & AESL_inst_dft.temp_94_loc_channel_U.if_full_n;
    assign fifo_intf_95.fifo_rd_block = 0;
    assign fifo_intf_95.fifo_wr_block = 0;
    assign fifo_intf_95.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_95;
    csv_file_dump cstatus_csv_dumper_95;
    df_fifo_monitor fifo_monitor_95;
    df_fifo_intf fifo_intf_96(clock,reset);
    assign fifo_intf_96.rd_en = AESL_inst_dft.temp_95_loc_channel_U.if_read & AESL_inst_dft.temp_95_loc_channel_U.if_empty_n;
    assign fifo_intf_96.wr_en = AESL_inst_dft.temp_95_loc_channel_U.if_write & AESL_inst_dft.temp_95_loc_channel_U.if_full_n;
    assign fifo_intf_96.fifo_rd_block = 0;
    assign fifo_intf_96.fifo_wr_block = 0;
    assign fifo_intf_96.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_96;
    csv_file_dump cstatus_csv_dumper_96;
    df_fifo_monitor fifo_monitor_96;
    df_fifo_intf fifo_intf_97(clock,reset);
    assign fifo_intf_97.rd_en = AESL_inst_dft.temp_96_loc_channel_U.if_read & AESL_inst_dft.temp_96_loc_channel_U.if_empty_n;
    assign fifo_intf_97.wr_en = AESL_inst_dft.temp_96_loc_channel_U.if_write & AESL_inst_dft.temp_96_loc_channel_U.if_full_n;
    assign fifo_intf_97.fifo_rd_block = 0;
    assign fifo_intf_97.fifo_wr_block = 0;
    assign fifo_intf_97.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_97;
    csv_file_dump cstatus_csv_dumper_97;
    df_fifo_monitor fifo_monitor_97;
    df_fifo_intf fifo_intf_98(clock,reset);
    assign fifo_intf_98.rd_en = AESL_inst_dft.temp_97_loc_channel_U.if_read & AESL_inst_dft.temp_97_loc_channel_U.if_empty_n;
    assign fifo_intf_98.wr_en = AESL_inst_dft.temp_97_loc_channel_U.if_write & AESL_inst_dft.temp_97_loc_channel_U.if_full_n;
    assign fifo_intf_98.fifo_rd_block = 0;
    assign fifo_intf_98.fifo_wr_block = 0;
    assign fifo_intf_98.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_98;
    csv_file_dump cstatus_csv_dumper_98;
    df_fifo_monitor fifo_monitor_98;
    df_fifo_intf fifo_intf_99(clock,reset);
    assign fifo_intf_99.rd_en = AESL_inst_dft.temp_98_loc_channel_U.if_read & AESL_inst_dft.temp_98_loc_channel_U.if_empty_n;
    assign fifo_intf_99.wr_en = AESL_inst_dft.temp_98_loc_channel_U.if_write & AESL_inst_dft.temp_98_loc_channel_U.if_full_n;
    assign fifo_intf_99.fifo_rd_block = 0;
    assign fifo_intf_99.fifo_wr_block = 0;
    assign fifo_intf_99.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_99;
    csv_file_dump cstatus_csv_dumper_99;
    df_fifo_monitor fifo_monitor_99;
    df_fifo_intf fifo_intf_100(clock,reset);
    assign fifo_intf_100.rd_en = AESL_inst_dft.temp_99_loc_channel_U.if_read & AESL_inst_dft.temp_99_loc_channel_U.if_empty_n;
    assign fifo_intf_100.wr_en = AESL_inst_dft.temp_99_loc_channel_U.if_write & AESL_inst_dft.temp_99_loc_channel_U.if_full_n;
    assign fifo_intf_100.fifo_rd_block = 0;
    assign fifo_intf_100.fifo_wr_block = 0;
    assign fifo_intf_100.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_100;
    csv_file_dump cstatus_csv_dumper_100;
    df_fifo_monitor fifo_monitor_100;
    df_fifo_intf fifo_intf_101(clock,reset);
    assign fifo_intf_101.rd_en = AESL_inst_dft.temp_100_loc_channel_U.if_read & AESL_inst_dft.temp_100_loc_channel_U.if_empty_n;
    assign fifo_intf_101.wr_en = AESL_inst_dft.temp_100_loc_channel_U.if_write & AESL_inst_dft.temp_100_loc_channel_U.if_full_n;
    assign fifo_intf_101.fifo_rd_block = 0;
    assign fifo_intf_101.fifo_wr_block = 0;
    assign fifo_intf_101.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_101;
    csv_file_dump cstatus_csv_dumper_101;
    df_fifo_monitor fifo_monitor_101;
    df_fifo_intf fifo_intf_102(clock,reset);
    assign fifo_intf_102.rd_en = AESL_inst_dft.temp_101_loc_channel_U.if_read & AESL_inst_dft.temp_101_loc_channel_U.if_empty_n;
    assign fifo_intf_102.wr_en = AESL_inst_dft.temp_101_loc_channel_U.if_write & AESL_inst_dft.temp_101_loc_channel_U.if_full_n;
    assign fifo_intf_102.fifo_rd_block = 0;
    assign fifo_intf_102.fifo_wr_block = 0;
    assign fifo_intf_102.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_102;
    csv_file_dump cstatus_csv_dumper_102;
    df_fifo_monitor fifo_monitor_102;
    df_fifo_intf fifo_intf_103(clock,reset);
    assign fifo_intf_103.rd_en = AESL_inst_dft.temp_102_loc_channel_U.if_read & AESL_inst_dft.temp_102_loc_channel_U.if_empty_n;
    assign fifo_intf_103.wr_en = AESL_inst_dft.temp_102_loc_channel_U.if_write & AESL_inst_dft.temp_102_loc_channel_U.if_full_n;
    assign fifo_intf_103.fifo_rd_block = 0;
    assign fifo_intf_103.fifo_wr_block = 0;
    assign fifo_intf_103.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_103;
    csv_file_dump cstatus_csv_dumper_103;
    df_fifo_monitor fifo_monitor_103;
    df_fifo_intf fifo_intf_104(clock,reset);
    assign fifo_intf_104.rd_en = AESL_inst_dft.temp_103_loc_channel_U.if_read & AESL_inst_dft.temp_103_loc_channel_U.if_empty_n;
    assign fifo_intf_104.wr_en = AESL_inst_dft.temp_103_loc_channel_U.if_write & AESL_inst_dft.temp_103_loc_channel_U.if_full_n;
    assign fifo_intf_104.fifo_rd_block = 0;
    assign fifo_intf_104.fifo_wr_block = 0;
    assign fifo_intf_104.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_104;
    csv_file_dump cstatus_csv_dumper_104;
    df_fifo_monitor fifo_monitor_104;
    df_fifo_intf fifo_intf_105(clock,reset);
    assign fifo_intf_105.rd_en = AESL_inst_dft.temp_104_loc_channel_U.if_read & AESL_inst_dft.temp_104_loc_channel_U.if_empty_n;
    assign fifo_intf_105.wr_en = AESL_inst_dft.temp_104_loc_channel_U.if_write & AESL_inst_dft.temp_104_loc_channel_U.if_full_n;
    assign fifo_intf_105.fifo_rd_block = 0;
    assign fifo_intf_105.fifo_wr_block = 0;
    assign fifo_intf_105.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_105;
    csv_file_dump cstatus_csv_dumper_105;
    df_fifo_monitor fifo_monitor_105;
    df_fifo_intf fifo_intf_106(clock,reset);
    assign fifo_intf_106.rd_en = AESL_inst_dft.temp_105_loc_channel_U.if_read & AESL_inst_dft.temp_105_loc_channel_U.if_empty_n;
    assign fifo_intf_106.wr_en = AESL_inst_dft.temp_105_loc_channel_U.if_write & AESL_inst_dft.temp_105_loc_channel_U.if_full_n;
    assign fifo_intf_106.fifo_rd_block = 0;
    assign fifo_intf_106.fifo_wr_block = 0;
    assign fifo_intf_106.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_106;
    csv_file_dump cstatus_csv_dumper_106;
    df_fifo_monitor fifo_monitor_106;
    df_fifo_intf fifo_intf_107(clock,reset);
    assign fifo_intf_107.rd_en = AESL_inst_dft.temp_106_loc_channel_U.if_read & AESL_inst_dft.temp_106_loc_channel_U.if_empty_n;
    assign fifo_intf_107.wr_en = AESL_inst_dft.temp_106_loc_channel_U.if_write & AESL_inst_dft.temp_106_loc_channel_U.if_full_n;
    assign fifo_intf_107.fifo_rd_block = 0;
    assign fifo_intf_107.fifo_wr_block = 0;
    assign fifo_intf_107.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_107;
    csv_file_dump cstatus_csv_dumper_107;
    df_fifo_monitor fifo_monitor_107;
    df_fifo_intf fifo_intf_108(clock,reset);
    assign fifo_intf_108.rd_en = AESL_inst_dft.temp_107_loc_channel_U.if_read & AESL_inst_dft.temp_107_loc_channel_U.if_empty_n;
    assign fifo_intf_108.wr_en = AESL_inst_dft.temp_107_loc_channel_U.if_write & AESL_inst_dft.temp_107_loc_channel_U.if_full_n;
    assign fifo_intf_108.fifo_rd_block = 0;
    assign fifo_intf_108.fifo_wr_block = 0;
    assign fifo_intf_108.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_108;
    csv_file_dump cstatus_csv_dumper_108;
    df_fifo_monitor fifo_monitor_108;
    df_fifo_intf fifo_intf_109(clock,reset);
    assign fifo_intf_109.rd_en = AESL_inst_dft.temp_108_loc_channel_U.if_read & AESL_inst_dft.temp_108_loc_channel_U.if_empty_n;
    assign fifo_intf_109.wr_en = AESL_inst_dft.temp_108_loc_channel_U.if_write & AESL_inst_dft.temp_108_loc_channel_U.if_full_n;
    assign fifo_intf_109.fifo_rd_block = 0;
    assign fifo_intf_109.fifo_wr_block = 0;
    assign fifo_intf_109.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_109;
    csv_file_dump cstatus_csv_dumper_109;
    df_fifo_monitor fifo_monitor_109;
    df_fifo_intf fifo_intf_110(clock,reset);
    assign fifo_intf_110.rd_en = AESL_inst_dft.temp_109_loc_channel_U.if_read & AESL_inst_dft.temp_109_loc_channel_U.if_empty_n;
    assign fifo_intf_110.wr_en = AESL_inst_dft.temp_109_loc_channel_U.if_write & AESL_inst_dft.temp_109_loc_channel_U.if_full_n;
    assign fifo_intf_110.fifo_rd_block = 0;
    assign fifo_intf_110.fifo_wr_block = 0;
    assign fifo_intf_110.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_110;
    csv_file_dump cstatus_csv_dumper_110;
    df_fifo_monitor fifo_monitor_110;
    df_fifo_intf fifo_intf_111(clock,reset);
    assign fifo_intf_111.rd_en = AESL_inst_dft.temp_110_loc_channel_U.if_read & AESL_inst_dft.temp_110_loc_channel_U.if_empty_n;
    assign fifo_intf_111.wr_en = AESL_inst_dft.temp_110_loc_channel_U.if_write & AESL_inst_dft.temp_110_loc_channel_U.if_full_n;
    assign fifo_intf_111.fifo_rd_block = 0;
    assign fifo_intf_111.fifo_wr_block = 0;
    assign fifo_intf_111.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_111;
    csv_file_dump cstatus_csv_dumper_111;
    df_fifo_monitor fifo_monitor_111;
    df_fifo_intf fifo_intf_112(clock,reset);
    assign fifo_intf_112.rd_en = AESL_inst_dft.temp_111_loc_channel_U.if_read & AESL_inst_dft.temp_111_loc_channel_U.if_empty_n;
    assign fifo_intf_112.wr_en = AESL_inst_dft.temp_111_loc_channel_U.if_write & AESL_inst_dft.temp_111_loc_channel_U.if_full_n;
    assign fifo_intf_112.fifo_rd_block = 0;
    assign fifo_intf_112.fifo_wr_block = 0;
    assign fifo_intf_112.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_112;
    csv_file_dump cstatus_csv_dumper_112;
    df_fifo_monitor fifo_monitor_112;
    df_fifo_intf fifo_intf_113(clock,reset);
    assign fifo_intf_113.rd_en = AESL_inst_dft.temp_112_loc_channel_U.if_read & AESL_inst_dft.temp_112_loc_channel_U.if_empty_n;
    assign fifo_intf_113.wr_en = AESL_inst_dft.temp_112_loc_channel_U.if_write & AESL_inst_dft.temp_112_loc_channel_U.if_full_n;
    assign fifo_intf_113.fifo_rd_block = 0;
    assign fifo_intf_113.fifo_wr_block = 0;
    assign fifo_intf_113.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_113;
    csv_file_dump cstatus_csv_dumper_113;
    df_fifo_monitor fifo_monitor_113;
    df_fifo_intf fifo_intf_114(clock,reset);
    assign fifo_intf_114.rd_en = AESL_inst_dft.temp_113_loc_channel_U.if_read & AESL_inst_dft.temp_113_loc_channel_U.if_empty_n;
    assign fifo_intf_114.wr_en = AESL_inst_dft.temp_113_loc_channel_U.if_write & AESL_inst_dft.temp_113_loc_channel_U.if_full_n;
    assign fifo_intf_114.fifo_rd_block = 0;
    assign fifo_intf_114.fifo_wr_block = 0;
    assign fifo_intf_114.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_114;
    csv_file_dump cstatus_csv_dumper_114;
    df_fifo_monitor fifo_monitor_114;
    df_fifo_intf fifo_intf_115(clock,reset);
    assign fifo_intf_115.rd_en = AESL_inst_dft.temp_114_loc_channel_U.if_read & AESL_inst_dft.temp_114_loc_channel_U.if_empty_n;
    assign fifo_intf_115.wr_en = AESL_inst_dft.temp_114_loc_channel_U.if_write & AESL_inst_dft.temp_114_loc_channel_U.if_full_n;
    assign fifo_intf_115.fifo_rd_block = 0;
    assign fifo_intf_115.fifo_wr_block = 0;
    assign fifo_intf_115.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_115;
    csv_file_dump cstatus_csv_dumper_115;
    df_fifo_monitor fifo_monitor_115;
    df_fifo_intf fifo_intf_116(clock,reset);
    assign fifo_intf_116.rd_en = AESL_inst_dft.temp_115_loc_channel_U.if_read & AESL_inst_dft.temp_115_loc_channel_U.if_empty_n;
    assign fifo_intf_116.wr_en = AESL_inst_dft.temp_115_loc_channel_U.if_write & AESL_inst_dft.temp_115_loc_channel_U.if_full_n;
    assign fifo_intf_116.fifo_rd_block = 0;
    assign fifo_intf_116.fifo_wr_block = 0;
    assign fifo_intf_116.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_116;
    csv_file_dump cstatus_csv_dumper_116;
    df_fifo_monitor fifo_monitor_116;
    df_fifo_intf fifo_intf_117(clock,reset);
    assign fifo_intf_117.rd_en = AESL_inst_dft.temp_116_loc_channel_U.if_read & AESL_inst_dft.temp_116_loc_channel_U.if_empty_n;
    assign fifo_intf_117.wr_en = AESL_inst_dft.temp_116_loc_channel_U.if_write & AESL_inst_dft.temp_116_loc_channel_U.if_full_n;
    assign fifo_intf_117.fifo_rd_block = 0;
    assign fifo_intf_117.fifo_wr_block = 0;
    assign fifo_intf_117.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_117;
    csv_file_dump cstatus_csv_dumper_117;
    df_fifo_monitor fifo_monitor_117;
    df_fifo_intf fifo_intf_118(clock,reset);
    assign fifo_intf_118.rd_en = AESL_inst_dft.temp_117_loc_channel_U.if_read & AESL_inst_dft.temp_117_loc_channel_U.if_empty_n;
    assign fifo_intf_118.wr_en = AESL_inst_dft.temp_117_loc_channel_U.if_write & AESL_inst_dft.temp_117_loc_channel_U.if_full_n;
    assign fifo_intf_118.fifo_rd_block = 0;
    assign fifo_intf_118.fifo_wr_block = 0;
    assign fifo_intf_118.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_118;
    csv_file_dump cstatus_csv_dumper_118;
    df_fifo_monitor fifo_monitor_118;
    df_fifo_intf fifo_intf_119(clock,reset);
    assign fifo_intf_119.rd_en = AESL_inst_dft.temp_118_loc_channel_U.if_read & AESL_inst_dft.temp_118_loc_channel_U.if_empty_n;
    assign fifo_intf_119.wr_en = AESL_inst_dft.temp_118_loc_channel_U.if_write & AESL_inst_dft.temp_118_loc_channel_U.if_full_n;
    assign fifo_intf_119.fifo_rd_block = 0;
    assign fifo_intf_119.fifo_wr_block = 0;
    assign fifo_intf_119.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_119;
    csv_file_dump cstatus_csv_dumper_119;
    df_fifo_monitor fifo_monitor_119;
    df_fifo_intf fifo_intf_120(clock,reset);
    assign fifo_intf_120.rd_en = AESL_inst_dft.temp_119_loc_channel_U.if_read & AESL_inst_dft.temp_119_loc_channel_U.if_empty_n;
    assign fifo_intf_120.wr_en = AESL_inst_dft.temp_119_loc_channel_U.if_write & AESL_inst_dft.temp_119_loc_channel_U.if_full_n;
    assign fifo_intf_120.fifo_rd_block = 0;
    assign fifo_intf_120.fifo_wr_block = 0;
    assign fifo_intf_120.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_120;
    csv_file_dump cstatus_csv_dumper_120;
    df_fifo_monitor fifo_monitor_120;
    df_fifo_intf fifo_intf_121(clock,reset);
    assign fifo_intf_121.rd_en = AESL_inst_dft.temp_120_loc_channel_U.if_read & AESL_inst_dft.temp_120_loc_channel_U.if_empty_n;
    assign fifo_intf_121.wr_en = AESL_inst_dft.temp_120_loc_channel_U.if_write & AESL_inst_dft.temp_120_loc_channel_U.if_full_n;
    assign fifo_intf_121.fifo_rd_block = 0;
    assign fifo_intf_121.fifo_wr_block = 0;
    assign fifo_intf_121.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_121;
    csv_file_dump cstatus_csv_dumper_121;
    df_fifo_monitor fifo_monitor_121;
    df_fifo_intf fifo_intf_122(clock,reset);
    assign fifo_intf_122.rd_en = AESL_inst_dft.temp_121_loc_channel_U.if_read & AESL_inst_dft.temp_121_loc_channel_U.if_empty_n;
    assign fifo_intf_122.wr_en = AESL_inst_dft.temp_121_loc_channel_U.if_write & AESL_inst_dft.temp_121_loc_channel_U.if_full_n;
    assign fifo_intf_122.fifo_rd_block = 0;
    assign fifo_intf_122.fifo_wr_block = 0;
    assign fifo_intf_122.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_122;
    csv_file_dump cstatus_csv_dumper_122;
    df_fifo_monitor fifo_monitor_122;
    df_fifo_intf fifo_intf_123(clock,reset);
    assign fifo_intf_123.rd_en = AESL_inst_dft.temp_122_loc_channel_U.if_read & AESL_inst_dft.temp_122_loc_channel_U.if_empty_n;
    assign fifo_intf_123.wr_en = AESL_inst_dft.temp_122_loc_channel_U.if_write & AESL_inst_dft.temp_122_loc_channel_U.if_full_n;
    assign fifo_intf_123.fifo_rd_block = 0;
    assign fifo_intf_123.fifo_wr_block = 0;
    assign fifo_intf_123.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_123;
    csv_file_dump cstatus_csv_dumper_123;
    df_fifo_monitor fifo_monitor_123;
    df_fifo_intf fifo_intf_124(clock,reset);
    assign fifo_intf_124.rd_en = AESL_inst_dft.temp_123_loc_channel_U.if_read & AESL_inst_dft.temp_123_loc_channel_U.if_empty_n;
    assign fifo_intf_124.wr_en = AESL_inst_dft.temp_123_loc_channel_U.if_write & AESL_inst_dft.temp_123_loc_channel_U.if_full_n;
    assign fifo_intf_124.fifo_rd_block = 0;
    assign fifo_intf_124.fifo_wr_block = 0;
    assign fifo_intf_124.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_124;
    csv_file_dump cstatus_csv_dumper_124;
    df_fifo_monitor fifo_monitor_124;
    df_fifo_intf fifo_intf_125(clock,reset);
    assign fifo_intf_125.rd_en = AESL_inst_dft.temp_124_loc_channel_U.if_read & AESL_inst_dft.temp_124_loc_channel_U.if_empty_n;
    assign fifo_intf_125.wr_en = AESL_inst_dft.temp_124_loc_channel_U.if_write & AESL_inst_dft.temp_124_loc_channel_U.if_full_n;
    assign fifo_intf_125.fifo_rd_block = 0;
    assign fifo_intf_125.fifo_wr_block = 0;
    assign fifo_intf_125.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_125;
    csv_file_dump cstatus_csv_dumper_125;
    df_fifo_monitor fifo_monitor_125;
    df_fifo_intf fifo_intf_126(clock,reset);
    assign fifo_intf_126.rd_en = AESL_inst_dft.temp_125_loc_channel_U.if_read & AESL_inst_dft.temp_125_loc_channel_U.if_empty_n;
    assign fifo_intf_126.wr_en = AESL_inst_dft.temp_125_loc_channel_U.if_write & AESL_inst_dft.temp_125_loc_channel_U.if_full_n;
    assign fifo_intf_126.fifo_rd_block = 0;
    assign fifo_intf_126.fifo_wr_block = 0;
    assign fifo_intf_126.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_126;
    csv_file_dump cstatus_csv_dumper_126;
    df_fifo_monitor fifo_monitor_126;
    df_fifo_intf fifo_intf_127(clock,reset);
    assign fifo_intf_127.rd_en = AESL_inst_dft.temp_126_loc_channel_U.if_read & AESL_inst_dft.temp_126_loc_channel_U.if_empty_n;
    assign fifo_intf_127.wr_en = AESL_inst_dft.temp_126_loc_channel_U.if_write & AESL_inst_dft.temp_126_loc_channel_U.if_full_n;
    assign fifo_intf_127.fifo_rd_block = 0;
    assign fifo_intf_127.fifo_wr_block = 0;
    assign fifo_intf_127.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_127;
    csv_file_dump cstatus_csv_dumper_127;
    df_fifo_monitor fifo_monitor_127;
    df_fifo_intf fifo_intf_128(clock,reset);
    assign fifo_intf_128.rd_en = AESL_inst_dft.temp_127_loc_channel_U.if_read & AESL_inst_dft.temp_127_loc_channel_U.if_empty_n;
    assign fifo_intf_128.wr_en = AESL_inst_dft.temp_127_loc_channel_U.if_write & AESL_inst_dft.temp_127_loc_channel_U.if_full_n;
    assign fifo_intf_128.fifo_rd_block = 0;
    assign fifo_intf_128.fifo_wr_block = 0;
    assign fifo_intf_128.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_128;
    csv_file_dump cstatus_csv_dumper_128;
    df_fifo_monitor fifo_monitor_128;
    df_fifo_intf fifo_intf_129(clock,reset);
    assign fifo_intf_129.rd_en = AESL_inst_dft.temp_128_loc_channel_U.if_read & AESL_inst_dft.temp_128_loc_channel_U.if_empty_n;
    assign fifo_intf_129.wr_en = AESL_inst_dft.temp_128_loc_channel_U.if_write & AESL_inst_dft.temp_128_loc_channel_U.if_full_n;
    assign fifo_intf_129.fifo_rd_block = 0;
    assign fifo_intf_129.fifo_wr_block = 0;
    assign fifo_intf_129.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_129;
    csv_file_dump cstatus_csv_dumper_129;
    df_fifo_monitor fifo_monitor_129;
    df_fifo_intf fifo_intf_130(clock,reset);
    assign fifo_intf_130.rd_en = AESL_inst_dft.temp_129_loc_channel_U.if_read & AESL_inst_dft.temp_129_loc_channel_U.if_empty_n;
    assign fifo_intf_130.wr_en = AESL_inst_dft.temp_129_loc_channel_U.if_write & AESL_inst_dft.temp_129_loc_channel_U.if_full_n;
    assign fifo_intf_130.fifo_rd_block = 0;
    assign fifo_intf_130.fifo_wr_block = 0;
    assign fifo_intf_130.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_130;
    csv_file_dump cstatus_csv_dumper_130;
    df_fifo_monitor fifo_monitor_130;
    df_fifo_intf fifo_intf_131(clock,reset);
    assign fifo_intf_131.rd_en = AESL_inst_dft.temp_130_loc_channel_U.if_read & AESL_inst_dft.temp_130_loc_channel_U.if_empty_n;
    assign fifo_intf_131.wr_en = AESL_inst_dft.temp_130_loc_channel_U.if_write & AESL_inst_dft.temp_130_loc_channel_U.if_full_n;
    assign fifo_intf_131.fifo_rd_block = 0;
    assign fifo_intf_131.fifo_wr_block = 0;
    assign fifo_intf_131.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_131;
    csv_file_dump cstatus_csv_dumper_131;
    df_fifo_monitor fifo_monitor_131;
    df_fifo_intf fifo_intf_132(clock,reset);
    assign fifo_intf_132.rd_en = AESL_inst_dft.temp_131_loc_channel_U.if_read & AESL_inst_dft.temp_131_loc_channel_U.if_empty_n;
    assign fifo_intf_132.wr_en = AESL_inst_dft.temp_131_loc_channel_U.if_write & AESL_inst_dft.temp_131_loc_channel_U.if_full_n;
    assign fifo_intf_132.fifo_rd_block = 0;
    assign fifo_intf_132.fifo_wr_block = 0;
    assign fifo_intf_132.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_132;
    csv_file_dump cstatus_csv_dumper_132;
    df_fifo_monitor fifo_monitor_132;
    df_fifo_intf fifo_intf_133(clock,reset);
    assign fifo_intf_133.rd_en = AESL_inst_dft.temp_132_loc_channel_U.if_read & AESL_inst_dft.temp_132_loc_channel_U.if_empty_n;
    assign fifo_intf_133.wr_en = AESL_inst_dft.temp_132_loc_channel_U.if_write & AESL_inst_dft.temp_132_loc_channel_U.if_full_n;
    assign fifo_intf_133.fifo_rd_block = 0;
    assign fifo_intf_133.fifo_wr_block = 0;
    assign fifo_intf_133.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_133;
    csv_file_dump cstatus_csv_dumper_133;
    df_fifo_monitor fifo_monitor_133;
    df_fifo_intf fifo_intf_134(clock,reset);
    assign fifo_intf_134.rd_en = AESL_inst_dft.temp_133_loc_channel_U.if_read & AESL_inst_dft.temp_133_loc_channel_U.if_empty_n;
    assign fifo_intf_134.wr_en = AESL_inst_dft.temp_133_loc_channel_U.if_write & AESL_inst_dft.temp_133_loc_channel_U.if_full_n;
    assign fifo_intf_134.fifo_rd_block = 0;
    assign fifo_intf_134.fifo_wr_block = 0;
    assign fifo_intf_134.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_134;
    csv_file_dump cstatus_csv_dumper_134;
    df_fifo_monitor fifo_monitor_134;
    df_fifo_intf fifo_intf_135(clock,reset);
    assign fifo_intf_135.rd_en = AESL_inst_dft.temp_134_loc_channel_U.if_read & AESL_inst_dft.temp_134_loc_channel_U.if_empty_n;
    assign fifo_intf_135.wr_en = AESL_inst_dft.temp_134_loc_channel_U.if_write & AESL_inst_dft.temp_134_loc_channel_U.if_full_n;
    assign fifo_intf_135.fifo_rd_block = 0;
    assign fifo_intf_135.fifo_wr_block = 0;
    assign fifo_intf_135.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_135;
    csv_file_dump cstatus_csv_dumper_135;
    df_fifo_monitor fifo_monitor_135;
    df_fifo_intf fifo_intf_136(clock,reset);
    assign fifo_intf_136.rd_en = AESL_inst_dft.temp_135_loc_channel_U.if_read & AESL_inst_dft.temp_135_loc_channel_U.if_empty_n;
    assign fifo_intf_136.wr_en = AESL_inst_dft.temp_135_loc_channel_U.if_write & AESL_inst_dft.temp_135_loc_channel_U.if_full_n;
    assign fifo_intf_136.fifo_rd_block = 0;
    assign fifo_intf_136.fifo_wr_block = 0;
    assign fifo_intf_136.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_136;
    csv_file_dump cstatus_csv_dumper_136;
    df_fifo_monitor fifo_monitor_136;
    df_fifo_intf fifo_intf_137(clock,reset);
    assign fifo_intf_137.rd_en = AESL_inst_dft.temp_136_loc_channel_U.if_read & AESL_inst_dft.temp_136_loc_channel_U.if_empty_n;
    assign fifo_intf_137.wr_en = AESL_inst_dft.temp_136_loc_channel_U.if_write & AESL_inst_dft.temp_136_loc_channel_U.if_full_n;
    assign fifo_intf_137.fifo_rd_block = 0;
    assign fifo_intf_137.fifo_wr_block = 0;
    assign fifo_intf_137.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_137;
    csv_file_dump cstatus_csv_dumper_137;
    df_fifo_monitor fifo_monitor_137;
    df_fifo_intf fifo_intf_138(clock,reset);
    assign fifo_intf_138.rd_en = AESL_inst_dft.temp_137_loc_channel_U.if_read & AESL_inst_dft.temp_137_loc_channel_U.if_empty_n;
    assign fifo_intf_138.wr_en = AESL_inst_dft.temp_137_loc_channel_U.if_write & AESL_inst_dft.temp_137_loc_channel_U.if_full_n;
    assign fifo_intf_138.fifo_rd_block = 0;
    assign fifo_intf_138.fifo_wr_block = 0;
    assign fifo_intf_138.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_138;
    csv_file_dump cstatus_csv_dumper_138;
    df_fifo_monitor fifo_monitor_138;
    df_fifo_intf fifo_intf_139(clock,reset);
    assign fifo_intf_139.rd_en = AESL_inst_dft.temp_138_loc_channel_U.if_read & AESL_inst_dft.temp_138_loc_channel_U.if_empty_n;
    assign fifo_intf_139.wr_en = AESL_inst_dft.temp_138_loc_channel_U.if_write & AESL_inst_dft.temp_138_loc_channel_U.if_full_n;
    assign fifo_intf_139.fifo_rd_block = 0;
    assign fifo_intf_139.fifo_wr_block = 0;
    assign fifo_intf_139.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_139;
    csv_file_dump cstatus_csv_dumper_139;
    df_fifo_monitor fifo_monitor_139;
    df_fifo_intf fifo_intf_140(clock,reset);
    assign fifo_intf_140.rd_en = AESL_inst_dft.temp_139_loc_channel_U.if_read & AESL_inst_dft.temp_139_loc_channel_U.if_empty_n;
    assign fifo_intf_140.wr_en = AESL_inst_dft.temp_139_loc_channel_U.if_write & AESL_inst_dft.temp_139_loc_channel_U.if_full_n;
    assign fifo_intf_140.fifo_rd_block = 0;
    assign fifo_intf_140.fifo_wr_block = 0;
    assign fifo_intf_140.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_140;
    csv_file_dump cstatus_csv_dumper_140;
    df_fifo_monitor fifo_monitor_140;
    df_fifo_intf fifo_intf_141(clock,reset);
    assign fifo_intf_141.rd_en = AESL_inst_dft.temp_140_loc_channel_U.if_read & AESL_inst_dft.temp_140_loc_channel_U.if_empty_n;
    assign fifo_intf_141.wr_en = AESL_inst_dft.temp_140_loc_channel_U.if_write & AESL_inst_dft.temp_140_loc_channel_U.if_full_n;
    assign fifo_intf_141.fifo_rd_block = 0;
    assign fifo_intf_141.fifo_wr_block = 0;
    assign fifo_intf_141.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_141;
    csv_file_dump cstatus_csv_dumper_141;
    df_fifo_monitor fifo_monitor_141;
    df_fifo_intf fifo_intf_142(clock,reset);
    assign fifo_intf_142.rd_en = AESL_inst_dft.temp_141_loc_channel_U.if_read & AESL_inst_dft.temp_141_loc_channel_U.if_empty_n;
    assign fifo_intf_142.wr_en = AESL_inst_dft.temp_141_loc_channel_U.if_write & AESL_inst_dft.temp_141_loc_channel_U.if_full_n;
    assign fifo_intf_142.fifo_rd_block = 0;
    assign fifo_intf_142.fifo_wr_block = 0;
    assign fifo_intf_142.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_142;
    csv_file_dump cstatus_csv_dumper_142;
    df_fifo_monitor fifo_monitor_142;
    df_fifo_intf fifo_intf_143(clock,reset);
    assign fifo_intf_143.rd_en = AESL_inst_dft.temp_142_loc_channel_U.if_read & AESL_inst_dft.temp_142_loc_channel_U.if_empty_n;
    assign fifo_intf_143.wr_en = AESL_inst_dft.temp_142_loc_channel_U.if_write & AESL_inst_dft.temp_142_loc_channel_U.if_full_n;
    assign fifo_intf_143.fifo_rd_block = 0;
    assign fifo_intf_143.fifo_wr_block = 0;
    assign fifo_intf_143.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_143;
    csv_file_dump cstatus_csv_dumper_143;
    df_fifo_monitor fifo_monitor_143;
    df_fifo_intf fifo_intf_144(clock,reset);
    assign fifo_intf_144.rd_en = AESL_inst_dft.temp_143_loc_channel_U.if_read & AESL_inst_dft.temp_143_loc_channel_U.if_empty_n;
    assign fifo_intf_144.wr_en = AESL_inst_dft.temp_143_loc_channel_U.if_write & AESL_inst_dft.temp_143_loc_channel_U.if_full_n;
    assign fifo_intf_144.fifo_rd_block = 0;
    assign fifo_intf_144.fifo_wr_block = 0;
    assign fifo_intf_144.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_144;
    csv_file_dump cstatus_csv_dumper_144;
    df_fifo_monitor fifo_monitor_144;
    df_fifo_intf fifo_intf_145(clock,reset);
    assign fifo_intf_145.rd_en = AESL_inst_dft.temp_144_loc_channel_U.if_read & AESL_inst_dft.temp_144_loc_channel_U.if_empty_n;
    assign fifo_intf_145.wr_en = AESL_inst_dft.temp_144_loc_channel_U.if_write & AESL_inst_dft.temp_144_loc_channel_U.if_full_n;
    assign fifo_intf_145.fifo_rd_block = 0;
    assign fifo_intf_145.fifo_wr_block = 0;
    assign fifo_intf_145.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_145;
    csv_file_dump cstatus_csv_dumper_145;
    df_fifo_monitor fifo_monitor_145;
    df_fifo_intf fifo_intf_146(clock,reset);
    assign fifo_intf_146.rd_en = AESL_inst_dft.temp_145_loc_channel_U.if_read & AESL_inst_dft.temp_145_loc_channel_U.if_empty_n;
    assign fifo_intf_146.wr_en = AESL_inst_dft.temp_145_loc_channel_U.if_write & AESL_inst_dft.temp_145_loc_channel_U.if_full_n;
    assign fifo_intf_146.fifo_rd_block = 0;
    assign fifo_intf_146.fifo_wr_block = 0;
    assign fifo_intf_146.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_146;
    csv_file_dump cstatus_csv_dumper_146;
    df_fifo_monitor fifo_monitor_146;
    df_fifo_intf fifo_intf_147(clock,reset);
    assign fifo_intf_147.rd_en = AESL_inst_dft.temp_146_loc_channel_U.if_read & AESL_inst_dft.temp_146_loc_channel_U.if_empty_n;
    assign fifo_intf_147.wr_en = AESL_inst_dft.temp_146_loc_channel_U.if_write & AESL_inst_dft.temp_146_loc_channel_U.if_full_n;
    assign fifo_intf_147.fifo_rd_block = 0;
    assign fifo_intf_147.fifo_wr_block = 0;
    assign fifo_intf_147.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_147;
    csv_file_dump cstatus_csv_dumper_147;
    df_fifo_monitor fifo_monitor_147;
    df_fifo_intf fifo_intf_148(clock,reset);
    assign fifo_intf_148.rd_en = AESL_inst_dft.temp_147_loc_channel_U.if_read & AESL_inst_dft.temp_147_loc_channel_U.if_empty_n;
    assign fifo_intf_148.wr_en = AESL_inst_dft.temp_147_loc_channel_U.if_write & AESL_inst_dft.temp_147_loc_channel_U.if_full_n;
    assign fifo_intf_148.fifo_rd_block = 0;
    assign fifo_intf_148.fifo_wr_block = 0;
    assign fifo_intf_148.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_148;
    csv_file_dump cstatus_csv_dumper_148;
    df_fifo_monitor fifo_monitor_148;
    df_fifo_intf fifo_intf_149(clock,reset);
    assign fifo_intf_149.rd_en = AESL_inst_dft.temp_148_loc_channel_U.if_read & AESL_inst_dft.temp_148_loc_channel_U.if_empty_n;
    assign fifo_intf_149.wr_en = AESL_inst_dft.temp_148_loc_channel_U.if_write & AESL_inst_dft.temp_148_loc_channel_U.if_full_n;
    assign fifo_intf_149.fifo_rd_block = 0;
    assign fifo_intf_149.fifo_wr_block = 0;
    assign fifo_intf_149.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_149;
    csv_file_dump cstatus_csv_dumper_149;
    df_fifo_monitor fifo_monitor_149;
    df_fifo_intf fifo_intf_150(clock,reset);
    assign fifo_intf_150.rd_en = AESL_inst_dft.temp_149_loc_channel_U.if_read & AESL_inst_dft.temp_149_loc_channel_U.if_empty_n;
    assign fifo_intf_150.wr_en = AESL_inst_dft.temp_149_loc_channel_U.if_write & AESL_inst_dft.temp_149_loc_channel_U.if_full_n;
    assign fifo_intf_150.fifo_rd_block = 0;
    assign fifo_intf_150.fifo_wr_block = 0;
    assign fifo_intf_150.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_150;
    csv_file_dump cstatus_csv_dumper_150;
    df_fifo_monitor fifo_monitor_150;
    df_fifo_intf fifo_intf_151(clock,reset);
    assign fifo_intf_151.rd_en = AESL_inst_dft.temp_150_loc_channel_U.if_read & AESL_inst_dft.temp_150_loc_channel_U.if_empty_n;
    assign fifo_intf_151.wr_en = AESL_inst_dft.temp_150_loc_channel_U.if_write & AESL_inst_dft.temp_150_loc_channel_U.if_full_n;
    assign fifo_intf_151.fifo_rd_block = 0;
    assign fifo_intf_151.fifo_wr_block = 0;
    assign fifo_intf_151.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_151;
    csv_file_dump cstatus_csv_dumper_151;
    df_fifo_monitor fifo_monitor_151;
    df_fifo_intf fifo_intf_152(clock,reset);
    assign fifo_intf_152.rd_en = AESL_inst_dft.temp_151_loc_channel_U.if_read & AESL_inst_dft.temp_151_loc_channel_U.if_empty_n;
    assign fifo_intf_152.wr_en = AESL_inst_dft.temp_151_loc_channel_U.if_write & AESL_inst_dft.temp_151_loc_channel_U.if_full_n;
    assign fifo_intf_152.fifo_rd_block = 0;
    assign fifo_intf_152.fifo_wr_block = 0;
    assign fifo_intf_152.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_152;
    csv_file_dump cstatus_csv_dumper_152;
    df_fifo_monitor fifo_monitor_152;
    df_fifo_intf fifo_intf_153(clock,reset);
    assign fifo_intf_153.rd_en = AESL_inst_dft.temp_152_loc_channel_U.if_read & AESL_inst_dft.temp_152_loc_channel_U.if_empty_n;
    assign fifo_intf_153.wr_en = AESL_inst_dft.temp_152_loc_channel_U.if_write & AESL_inst_dft.temp_152_loc_channel_U.if_full_n;
    assign fifo_intf_153.fifo_rd_block = 0;
    assign fifo_intf_153.fifo_wr_block = 0;
    assign fifo_intf_153.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_153;
    csv_file_dump cstatus_csv_dumper_153;
    df_fifo_monitor fifo_monitor_153;
    df_fifo_intf fifo_intf_154(clock,reset);
    assign fifo_intf_154.rd_en = AESL_inst_dft.temp_153_loc_channel_U.if_read & AESL_inst_dft.temp_153_loc_channel_U.if_empty_n;
    assign fifo_intf_154.wr_en = AESL_inst_dft.temp_153_loc_channel_U.if_write & AESL_inst_dft.temp_153_loc_channel_U.if_full_n;
    assign fifo_intf_154.fifo_rd_block = 0;
    assign fifo_intf_154.fifo_wr_block = 0;
    assign fifo_intf_154.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_154;
    csv_file_dump cstatus_csv_dumper_154;
    df_fifo_monitor fifo_monitor_154;
    df_fifo_intf fifo_intf_155(clock,reset);
    assign fifo_intf_155.rd_en = AESL_inst_dft.temp_154_loc_channel_U.if_read & AESL_inst_dft.temp_154_loc_channel_U.if_empty_n;
    assign fifo_intf_155.wr_en = AESL_inst_dft.temp_154_loc_channel_U.if_write & AESL_inst_dft.temp_154_loc_channel_U.if_full_n;
    assign fifo_intf_155.fifo_rd_block = 0;
    assign fifo_intf_155.fifo_wr_block = 0;
    assign fifo_intf_155.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_155;
    csv_file_dump cstatus_csv_dumper_155;
    df_fifo_monitor fifo_monitor_155;
    df_fifo_intf fifo_intf_156(clock,reset);
    assign fifo_intf_156.rd_en = AESL_inst_dft.temp_155_loc_channel_U.if_read & AESL_inst_dft.temp_155_loc_channel_U.if_empty_n;
    assign fifo_intf_156.wr_en = AESL_inst_dft.temp_155_loc_channel_U.if_write & AESL_inst_dft.temp_155_loc_channel_U.if_full_n;
    assign fifo_intf_156.fifo_rd_block = 0;
    assign fifo_intf_156.fifo_wr_block = 0;
    assign fifo_intf_156.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_156;
    csv_file_dump cstatus_csv_dumper_156;
    df_fifo_monitor fifo_monitor_156;
    df_fifo_intf fifo_intf_157(clock,reset);
    assign fifo_intf_157.rd_en = AESL_inst_dft.temp_156_loc_channel_U.if_read & AESL_inst_dft.temp_156_loc_channel_U.if_empty_n;
    assign fifo_intf_157.wr_en = AESL_inst_dft.temp_156_loc_channel_U.if_write & AESL_inst_dft.temp_156_loc_channel_U.if_full_n;
    assign fifo_intf_157.fifo_rd_block = 0;
    assign fifo_intf_157.fifo_wr_block = 0;
    assign fifo_intf_157.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_157;
    csv_file_dump cstatus_csv_dumper_157;
    df_fifo_monitor fifo_monitor_157;
    df_fifo_intf fifo_intf_158(clock,reset);
    assign fifo_intf_158.rd_en = AESL_inst_dft.temp_157_loc_channel_U.if_read & AESL_inst_dft.temp_157_loc_channel_U.if_empty_n;
    assign fifo_intf_158.wr_en = AESL_inst_dft.temp_157_loc_channel_U.if_write & AESL_inst_dft.temp_157_loc_channel_U.if_full_n;
    assign fifo_intf_158.fifo_rd_block = 0;
    assign fifo_intf_158.fifo_wr_block = 0;
    assign fifo_intf_158.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_158;
    csv_file_dump cstatus_csv_dumper_158;
    df_fifo_monitor fifo_monitor_158;
    df_fifo_intf fifo_intf_159(clock,reset);
    assign fifo_intf_159.rd_en = AESL_inst_dft.temp_158_loc_channel_U.if_read & AESL_inst_dft.temp_158_loc_channel_U.if_empty_n;
    assign fifo_intf_159.wr_en = AESL_inst_dft.temp_158_loc_channel_U.if_write & AESL_inst_dft.temp_158_loc_channel_U.if_full_n;
    assign fifo_intf_159.fifo_rd_block = 0;
    assign fifo_intf_159.fifo_wr_block = 0;
    assign fifo_intf_159.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_159;
    csv_file_dump cstatus_csv_dumper_159;
    df_fifo_monitor fifo_monitor_159;
    df_fifo_intf fifo_intf_160(clock,reset);
    assign fifo_intf_160.rd_en = AESL_inst_dft.temp_159_loc_channel_U.if_read & AESL_inst_dft.temp_159_loc_channel_U.if_empty_n;
    assign fifo_intf_160.wr_en = AESL_inst_dft.temp_159_loc_channel_U.if_write & AESL_inst_dft.temp_159_loc_channel_U.if_full_n;
    assign fifo_intf_160.fifo_rd_block = 0;
    assign fifo_intf_160.fifo_wr_block = 0;
    assign fifo_intf_160.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_160;
    csv_file_dump cstatus_csv_dumper_160;
    df_fifo_monitor fifo_monitor_160;
    df_fifo_intf fifo_intf_161(clock,reset);
    assign fifo_intf_161.rd_en = AESL_inst_dft.temp_160_loc_channel_U.if_read & AESL_inst_dft.temp_160_loc_channel_U.if_empty_n;
    assign fifo_intf_161.wr_en = AESL_inst_dft.temp_160_loc_channel_U.if_write & AESL_inst_dft.temp_160_loc_channel_U.if_full_n;
    assign fifo_intf_161.fifo_rd_block = 0;
    assign fifo_intf_161.fifo_wr_block = 0;
    assign fifo_intf_161.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_161;
    csv_file_dump cstatus_csv_dumper_161;
    df_fifo_monitor fifo_monitor_161;
    df_fifo_intf fifo_intf_162(clock,reset);
    assign fifo_intf_162.rd_en = AESL_inst_dft.temp_161_loc_channel_U.if_read & AESL_inst_dft.temp_161_loc_channel_U.if_empty_n;
    assign fifo_intf_162.wr_en = AESL_inst_dft.temp_161_loc_channel_U.if_write & AESL_inst_dft.temp_161_loc_channel_U.if_full_n;
    assign fifo_intf_162.fifo_rd_block = 0;
    assign fifo_intf_162.fifo_wr_block = 0;
    assign fifo_intf_162.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_162;
    csv_file_dump cstatus_csv_dumper_162;
    df_fifo_monitor fifo_monitor_162;
    df_fifo_intf fifo_intf_163(clock,reset);
    assign fifo_intf_163.rd_en = AESL_inst_dft.temp_162_loc_channel_U.if_read & AESL_inst_dft.temp_162_loc_channel_U.if_empty_n;
    assign fifo_intf_163.wr_en = AESL_inst_dft.temp_162_loc_channel_U.if_write & AESL_inst_dft.temp_162_loc_channel_U.if_full_n;
    assign fifo_intf_163.fifo_rd_block = 0;
    assign fifo_intf_163.fifo_wr_block = 0;
    assign fifo_intf_163.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_163;
    csv_file_dump cstatus_csv_dumper_163;
    df_fifo_monitor fifo_monitor_163;
    df_fifo_intf fifo_intf_164(clock,reset);
    assign fifo_intf_164.rd_en = AESL_inst_dft.temp_163_loc_channel_U.if_read & AESL_inst_dft.temp_163_loc_channel_U.if_empty_n;
    assign fifo_intf_164.wr_en = AESL_inst_dft.temp_163_loc_channel_U.if_write & AESL_inst_dft.temp_163_loc_channel_U.if_full_n;
    assign fifo_intf_164.fifo_rd_block = 0;
    assign fifo_intf_164.fifo_wr_block = 0;
    assign fifo_intf_164.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_164;
    csv_file_dump cstatus_csv_dumper_164;
    df_fifo_monitor fifo_monitor_164;
    df_fifo_intf fifo_intf_165(clock,reset);
    assign fifo_intf_165.rd_en = AESL_inst_dft.temp_164_loc_channel_U.if_read & AESL_inst_dft.temp_164_loc_channel_U.if_empty_n;
    assign fifo_intf_165.wr_en = AESL_inst_dft.temp_164_loc_channel_U.if_write & AESL_inst_dft.temp_164_loc_channel_U.if_full_n;
    assign fifo_intf_165.fifo_rd_block = 0;
    assign fifo_intf_165.fifo_wr_block = 0;
    assign fifo_intf_165.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_165;
    csv_file_dump cstatus_csv_dumper_165;
    df_fifo_monitor fifo_monitor_165;
    df_fifo_intf fifo_intf_166(clock,reset);
    assign fifo_intf_166.rd_en = AESL_inst_dft.temp_165_loc_channel_U.if_read & AESL_inst_dft.temp_165_loc_channel_U.if_empty_n;
    assign fifo_intf_166.wr_en = AESL_inst_dft.temp_165_loc_channel_U.if_write & AESL_inst_dft.temp_165_loc_channel_U.if_full_n;
    assign fifo_intf_166.fifo_rd_block = 0;
    assign fifo_intf_166.fifo_wr_block = 0;
    assign fifo_intf_166.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_166;
    csv_file_dump cstatus_csv_dumper_166;
    df_fifo_monitor fifo_monitor_166;
    df_fifo_intf fifo_intf_167(clock,reset);
    assign fifo_intf_167.rd_en = AESL_inst_dft.temp_166_loc_channel_U.if_read & AESL_inst_dft.temp_166_loc_channel_U.if_empty_n;
    assign fifo_intf_167.wr_en = AESL_inst_dft.temp_166_loc_channel_U.if_write & AESL_inst_dft.temp_166_loc_channel_U.if_full_n;
    assign fifo_intf_167.fifo_rd_block = 0;
    assign fifo_intf_167.fifo_wr_block = 0;
    assign fifo_intf_167.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_167;
    csv_file_dump cstatus_csv_dumper_167;
    df_fifo_monitor fifo_monitor_167;
    df_fifo_intf fifo_intf_168(clock,reset);
    assign fifo_intf_168.rd_en = AESL_inst_dft.temp_167_loc_channel_U.if_read & AESL_inst_dft.temp_167_loc_channel_U.if_empty_n;
    assign fifo_intf_168.wr_en = AESL_inst_dft.temp_167_loc_channel_U.if_write & AESL_inst_dft.temp_167_loc_channel_U.if_full_n;
    assign fifo_intf_168.fifo_rd_block = 0;
    assign fifo_intf_168.fifo_wr_block = 0;
    assign fifo_intf_168.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_168;
    csv_file_dump cstatus_csv_dumper_168;
    df_fifo_monitor fifo_monitor_168;
    df_fifo_intf fifo_intf_169(clock,reset);
    assign fifo_intf_169.rd_en = AESL_inst_dft.temp_168_loc_channel_U.if_read & AESL_inst_dft.temp_168_loc_channel_U.if_empty_n;
    assign fifo_intf_169.wr_en = AESL_inst_dft.temp_168_loc_channel_U.if_write & AESL_inst_dft.temp_168_loc_channel_U.if_full_n;
    assign fifo_intf_169.fifo_rd_block = 0;
    assign fifo_intf_169.fifo_wr_block = 0;
    assign fifo_intf_169.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_169;
    csv_file_dump cstatus_csv_dumper_169;
    df_fifo_monitor fifo_monitor_169;
    df_fifo_intf fifo_intf_170(clock,reset);
    assign fifo_intf_170.rd_en = AESL_inst_dft.temp_169_loc_channel_U.if_read & AESL_inst_dft.temp_169_loc_channel_U.if_empty_n;
    assign fifo_intf_170.wr_en = AESL_inst_dft.temp_169_loc_channel_U.if_write & AESL_inst_dft.temp_169_loc_channel_U.if_full_n;
    assign fifo_intf_170.fifo_rd_block = 0;
    assign fifo_intf_170.fifo_wr_block = 0;
    assign fifo_intf_170.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_170;
    csv_file_dump cstatus_csv_dumper_170;
    df_fifo_monitor fifo_monitor_170;
    df_fifo_intf fifo_intf_171(clock,reset);
    assign fifo_intf_171.rd_en = AESL_inst_dft.temp_170_loc_channel_U.if_read & AESL_inst_dft.temp_170_loc_channel_U.if_empty_n;
    assign fifo_intf_171.wr_en = AESL_inst_dft.temp_170_loc_channel_U.if_write & AESL_inst_dft.temp_170_loc_channel_U.if_full_n;
    assign fifo_intf_171.fifo_rd_block = 0;
    assign fifo_intf_171.fifo_wr_block = 0;
    assign fifo_intf_171.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_171;
    csv_file_dump cstatus_csv_dumper_171;
    df_fifo_monitor fifo_monitor_171;
    df_fifo_intf fifo_intf_172(clock,reset);
    assign fifo_intf_172.rd_en = AESL_inst_dft.temp_171_loc_channel_U.if_read & AESL_inst_dft.temp_171_loc_channel_U.if_empty_n;
    assign fifo_intf_172.wr_en = AESL_inst_dft.temp_171_loc_channel_U.if_write & AESL_inst_dft.temp_171_loc_channel_U.if_full_n;
    assign fifo_intf_172.fifo_rd_block = 0;
    assign fifo_intf_172.fifo_wr_block = 0;
    assign fifo_intf_172.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_172;
    csv_file_dump cstatus_csv_dumper_172;
    df_fifo_monitor fifo_monitor_172;
    df_fifo_intf fifo_intf_173(clock,reset);
    assign fifo_intf_173.rd_en = AESL_inst_dft.temp_172_loc_channel_U.if_read & AESL_inst_dft.temp_172_loc_channel_U.if_empty_n;
    assign fifo_intf_173.wr_en = AESL_inst_dft.temp_172_loc_channel_U.if_write & AESL_inst_dft.temp_172_loc_channel_U.if_full_n;
    assign fifo_intf_173.fifo_rd_block = 0;
    assign fifo_intf_173.fifo_wr_block = 0;
    assign fifo_intf_173.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_173;
    csv_file_dump cstatus_csv_dumper_173;
    df_fifo_monitor fifo_monitor_173;
    df_fifo_intf fifo_intf_174(clock,reset);
    assign fifo_intf_174.rd_en = AESL_inst_dft.temp_173_loc_channel_U.if_read & AESL_inst_dft.temp_173_loc_channel_U.if_empty_n;
    assign fifo_intf_174.wr_en = AESL_inst_dft.temp_173_loc_channel_U.if_write & AESL_inst_dft.temp_173_loc_channel_U.if_full_n;
    assign fifo_intf_174.fifo_rd_block = 0;
    assign fifo_intf_174.fifo_wr_block = 0;
    assign fifo_intf_174.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_174;
    csv_file_dump cstatus_csv_dumper_174;
    df_fifo_monitor fifo_monitor_174;
    df_fifo_intf fifo_intf_175(clock,reset);
    assign fifo_intf_175.rd_en = AESL_inst_dft.temp_174_loc_channel_U.if_read & AESL_inst_dft.temp_174_loc_channel_U.if_empty_n;
    assign fifo_intf_175.wr_en = AESL_inst_dft.temp_174_loc_channel_U.if_write & AESL_inst_dft.temp_174_loc_channel_U.if_full_n;
    assign fifo_intf_175.fifo_rd_block = 0;
    assign fifo_intf_175.fifo_wr_block = 0;
    assign fifo_intf_175.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_175;
    csv_file_dump cstatus_csv_dumper_175;
    df_fifo_monitor fifo_monitor_175;
    df_fifo_intf fifo_intf_176(clock,reset);
    assign fifo_intf_176.rd_en = AESL_inst_dft.temp_175_loc_channel_U.if_read & AESL_inst_dft.temp_175_loc_channel_U.if_empty_n;
    assign fifo_intf_176.wr_en = AESL_inst_dft.temp_175_loc_channel_U.if_write & AESL_inst_dft.temp_175_loc_channel_U.if_full_n;
    assign fifo_intf_176.fifo_rd_block = 0;
    assign fifo_intf_176.fifo_wr_block = 0;
    assign fifo_intf_176.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_176;
    csv_file_dump cstatus_csv_dumper_176;
    df_fifo_monitor fifo_monitor_176;
    df_fifo_intf fifo_intf_177(clock,reset);
    assign fifo_intf_177.rd_en = AESL_inst_dft.temp_176_loc_channel_U.if_read & AESL_inst_dft.temp_176_loc_channel_U.if_empty_n;
    assign fifo_intf_177.wr_en = AESL_inst_dft.temp_176_loc_channel_U.if_write & AESL_inst_dft.temp_176_loc_channel_U.if_full_n;
    assign fifo_intf_177.fifo_rd_block = 0;
    assign fifo_intf_177.fifo_wr_block = 0;
    assign fifo_intf_177.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_177;
    csv_file_dump cstatus_csv_dumper_177;
    df_fifo_monitor fifo_monitor_177;
    df_fifo_intf fifo_intf_178(clock,reset);
    assign fifo_intf_178.rd_en = AESL_inst_dft.temp_177_loc_channel_U.if_read & AESL_inst_dft.temp_177_loc_channel_U.if_empty_n;
    assign fifo_intf_178.wr_en = AESL_inst_dft.temp_177_loc_channel_U.if_write & AESL_inst_dft.temp_177_loc_channel_U.if_full_n;
    assign fifo_intf_178.fifo_rd_block = 0;
    assign fifo_intf_178.fifo_wr_block = 0;
    assign fifo_intf_178.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_178;
    csv_file_dump cstatus_csv_dumper_178;
    df_fifo_monitor fifo_monitor_178;
    df_fifo_intf fifo_intf_179(clock,reset);
    assign fifo_intf_179.rd_en = AESL_inst_dft.temp_178_loc_channel_U.if_read & AESL_inst_dft.temp_178_loc_channel_U.if_empty_n;
    assign fifo_intf_179.wr_en = AESL_inst_dft.temp_178_loc_channel_U.if_write & AESL_inst_dft.temp_178_loc_channel_U.if_full_n;
    assign fifo_intf_179.fifo_rd_block = 0;
    assign fifo_intf_179.fifo_wr_block = 0;
    assign fifo_intf_179.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_179;
    csv_file_dump cstatus_csv_dumper_179;
    df_fifo_monitor fifo_monitor_179;
    df_fifo_intf fifo_intf_180(clock,reset);
    assign fifo_intf_180.rd_en = AESL_inst_dft.temp_179_loc_channel_U.if_read & AESL_inst_dft.temp_179_loc_channel_U.if_empty_n;
    assign fifo_intf_180.wr_en = AESL_inst_dft.temp_179_loc_channel_U.if_write & AESL_inst_dft.temp_179_loc_channel_U.if_full_n;
    assign fifo_intf_180.fifo_rd_block = 0;
    assign fifo_intf_180.fifo_wr_block = 0;
    assign fifo_intf_180.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_180;
    csv_file_dump cstatus_csv_dumper_180;
    df_fifo_monitor fifo_monitor_180;
    df_fifo_intf fifo_intf_181(clock,reset);
    assign fifo_intf_181.rd_en = AESL_inst_dft.temp_180_loc_channel_U.if_read & AESL_inst_dft.temp_180_loc_channel_U.if_empty_n;
    assign fifo_intf_181.wr_en = AESL_inst_dft.temp_180_loc_channel_U.if_write & AESL_inst_dft.temp_180_loc_channel_U.if_full_n;
    assign fifo_intf_181.fifo_rd_block = 0;
    assign fifo_intf_181.fifo_wr_block = 0;
    assign fifo_intf_181.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_181;
    csv_file_dump cstatus_csv_dumper_181;
    df_fifo_monitor fifo_monitor_181;
    df_fifo_intf fifo_intf_182(clock,reset);
    assign fifo_intf_182.rd_en = AESL_inst_dft.temp_181_loc_channel_U.if_read & AESL_inst_dft.temp_181_loc_channel_U.if_empty_n;
    assign fifo_intf_182.wr_en = AESL_inst_dft.temp_181_loc_channel_U.if_write & AESL_inst_dft.temp_181_loc_channel_U.if_full_n;
    assign fifo_intf_182.fifo_rd_block = 0;
    assign fifo_intf_182.fifo_wr_block = 0;
    assign fifo_intf_182.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_182;
    csv_file_dump cstatus_csv_dumper_182;
    df_fifo_monitor fifo_monitor_182;
    df_fifo_intf fifo_intf_183(clock,reset);
    assign fifo_intf_183.rd_en = AESL_inst_dft.temp_182_loc_channel_U.if_read & AESL_inst_dft.temp_182_loc_channel_U.if_empty_n;
    assign fifo_intf_183.wr_en = AESL_inst_dft.temp_182_loc_channel_U.if_write & AESL_inst_dft.temp_182_loc_channel_U.if_full_n;
    assign fifo_intf_183.fifo_rd_block = 0;
    assign fifo_intf_183.fifo_wr_block = 0;
    assign fifo_intf_183.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_183;
    csv_file_dump cstatus_csv_dumper_183;
    df_fifo_monitor fifo_monitor_183;
    df_fifo_intf fifo_intf_184(clock,reset);
    assign fifo_intf_184.rd_en = AESL_inst_dft.temp_183_loc_channel_U.if_read & AESL_inst_dft.temp_183_loc_channel_U.if_empty_n;
    assign fifo_intf_184.wr_en = AESL_inst_dft.temp_183_loc_channel_U.if_write & AESL_inst_dft.temp_183_loc_channel_U.if_full_n;
    assign fifo_intf_184.fifo_rd_block = 0;
    assign fifo_intf_184.fifo_wr_block = 0;
    assign fifo_intf_184.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_184;
    csv_file_dump cstatus_csv_dumper_184;
    df_fifo_monitor fifo_monitor_184;
    df_fifo_intf fifo_intf_185(clock,reset);
    assign fifo_intf_185.rd_en = AESL_inst_dft.temp_184_loc_channel_U.if_read & AESL_inst_dft.temp_184_loc_channel_U.if_empty_n;
    assign fifo_intf_185.wr_en = AESL_inst_dft.temp_184_loc_channel_U.if_write & AESL_inst_dft.temp_184_loc_channel_U.if_full_n;
    assign fifo_intf_185.fifo_rd_block = 0;
    assign fifo_intf_185.fifo_wr_block = 0;
    assign fifo_intf_185.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_185;
    csv_file_dump cstatus_csv_dumper_185;
    df_fifo_monitor fifo_monitor_185;
    df_fifo_intf fifo_intf_186(clock,reset);
    assign fifo_intf_186.rd_en = AESL_inst_dft.temp_185_loc_channel_U.if_read & AESL_inst_dft.temp_185_loc_channel_U.if_empty_n;
    assign fifo_intf_186.wr_en = AESL_inst_dft.temp_185_loc_channel_U.if_write & AESL_inst_dft.temp_185_loc_channel_U.if_full_n;
    assign fifo_intf_186.fifo_rd_block = 0;
    assign fifo_intf_186.fifo_wr_block = 0;
    assign fifo_intf_186.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_186;
    csv_file_dump cstatus_csv_dumper_186;
    df_fifo_monitor fifo_monitor_186;
    df_fifo_intf fifo_intf_187(clock,reset);
    assign fifo_intf_187.rd_en = AESL_inst_dft.temp_186_loc_channel_U.if_read & AESL_inst_dft.temp_186_loc_channel_U.if_empty_n;
    assign fifo_intf_187.wr_en = AESL_inst_dft.temp_186_loc_channel_U.if_write & AESL_inst_dft.temp_186_loc_channel_U.if_full_n;
    assign fifo_intf_187.fifo_rd_block = 0;
    assign fifo_intf_187.fifo_wr_block = 0;
    assign fifo_intf_187.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_187;
    csv_file_dump cstatus_csv_dumper_187;
    df_fifo_monitor fifo_monitor_187;
    df_fifo_intf fifo_intf_188(clock,reset);
    assign fifo_intf_188.rd_en = AESL_inst_dft.temp_187_loc_channel_U.if_read & AESL_inst_dft.temp_187_loc_channel_U.if_empty_n;
    assign fifo_intf_188.wr_en = AESL_inst_dft.temp_187_loc_channel_U.if_write & AESL_inst_dft.temp_187_loc_channel_U.if_full_n;
    assign fifo_intf_188.fifo_rd_block = 0;
    assign fifo_intf_188.fifo_wr_block = 0;
    assign fifo_intf_188.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_188;
    csv_file_dump cstatus_csv_dumper_188;
    df_fifo_monitor fifo_monitor_188;
    df_fifo_intf fifo_intf_189(clock,reset);
    assign fifo_intf_189.rd_en = AESL_inst_dft.temp_188_loc_channel_U.if_read & AESL_inst_dft.temp_188_loc_channel_U.if_empty_n;
    assign fifo_intf_189.wr_en = AESL_inst_dft.temp_188_loc_channel_U.if_write & AESL_inst_dft.temp_188_loc_channel_U.if_full_n;
    assign fifo_intf_189.fifo_rd_block = 0;
    assign fifo_intf_189.fifo_wr_block = 0;
    assign fifo_intf_189.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_189;
    csv_file_dump cstatus_csv_dumper_189;
    df_fifo_monitor fifo_monitor_189;
    df_fifo_intf fifo_intf_190(clock,reset);
    assign fifo_intf_190.rd_en = AESL_inst_dft.temp_189_loc_channel_U.if_read & AESL_inst_dft.temp_189_loc_channel_U.if_empty_n;
    assign fifo_intf_190.wr_en = AESL_inst_dft.temp_189_loc_channel_U.if_write & AESL_inst_dft.temp_189_loc_channel_U.if_full_n;
    assign fifo_intf_190.fifo_rd_block = 0;
    assign fifo_intf_190.fifo_wr_block = 0;
    assign fifo_intf_190.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_190;
    csv_file_dump cstatus_csv_dumper_190;
    df_fifo_monitor fifo_monitor_190;
    df_fifo_intf fifo_intf_191(clock,reset);
    assign fifo_intf_191.rd_en = AESL_inst_dft.temp_190_loc_channel_U.if_read & AESL_inst_dft.temp_190_loc_channel_U.if_empty_n;
    assign fifo_intf_191.wr_en = AESL_inst_dft.temp_190_loc_channel_U.if_write & AESL_inst_dft.temp_190_loc_channel_U.if_full_n;
    assign fifo_intf_191.fifo_rd_block = 0;
    assign fifo_intf_191.fifo_wr_block = 0;
    assign fifo_intf_191.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_191;
    csv_file_dump cstatus_csv_dumper_191;
    df_fifo_monitor fifo_monitor_191;
    df_fifo_intf fifo_intf_192(clock,reset);
    assign fifo_intf_192.rd_en = AESL_inst_dft.temp_191_loc_channel_U.if_read & AESL_inst_dft.temp_191_loc_channel_U.if_empty_n;
    assign fifo_intf_192.wr_en = AESL_inst_dft.temp_191_loc_channel_U.if_write & AESL_inst_dft.temp_191_loc_channel_U.if_full_n;
    assign fifo_intf_192.fifo_rd_block = 0;
    assign fifo_intf_192.fifo_wr_block = 0;
    assign fifo_intf_192.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_192;
    csv_file_dump cstatus_csv_dumper_192;
    df_fifo_monitor fifo_monitor_192;
    df_fifo_intf fifo_intf_193(clock,reset);
    assign fifo_intf_193.rd_en = AESL_inst_dft.temp_192_loc_channel_U.if_read & AESL_inst_dft.temp_192_loc_channel_U.if_empty_n;
    assign fifo_intf_193.wr_en = AESL_inst_dft.temp_192_loc_channel_U.if_write & AESL_inst_dft.temp_192_loc_channel_U.if_full_n;
    assign fifo_intf_193.fifo_rd_block = 0;
    assign fifo_intf_193.fifo_wr_block = 0;
    assign fifo_intf_193.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_193;
    csv_file_dump cstatus_csv_dumper_193;
    df_fifo_monitor fifo_monitor_193;
    df_fifo_intf fifo_intf_194(clock,reset);
    assign fifo_intf_194.rd_en = AESL_inst_dft.temp_193_loc_channel_U.if_read & AESL_inst_dft.temp_193_loc_channel_U.if_empty_n;
    assign fifo_intf_194.wr_en = AESL_inst_dft.temp_193_loc_channel_U.if_write & AESL_inst_dft.temp_193_loc_channel_U.if_full_n;
    assign fifo_intf_194.fifo_rd_block = 0;
    assign fifo_intf_194.fifo_wr_block = 0;
    assign fifo_intf_194.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_194;
    csv_file_dump cstatus_csv_dumper_194;
    df_fifo_monitor fifo_monitor_194;
    df_fifo_intf fifo_intf_195(clock,reset);
    assign fifo_intf_195.rd_en = AESL_inst_dft.temp_194_loc_channel_U.if_read & AESL_inst_dft.temp_194_loc_channel_U.if_empty_n;
    assign fifo_intf_195.wr_en = AESL_inst_dft.temp_194_loc_channel_U.if_write & AESL_inst_dft.temp_194_loc_channel_U.if_full_n;
    assign fifo_intf_195.fifo_rd_block = 0;
    assign fifo_intf_195.fifo_wr_block = 0;
    assign fifo_intf_195.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_195;
    csv_file_dump cstatus_csv_dumper_195;
    df_fifo_monitor fifo_monitor_195;
    df_fifo_intf fifo_intf_196(clock,reset);
    assign fifo_intf_196.rd_en = AESL_inst_dft.temp_195_loc_channel_U.if_read & AESL_inst_dft.temp_195_loc_channel_U.if_empty_n;
    assign fifo_intf_196.wr_en = AESL_inst_dft.temp_195_loc_channel_U.if_write & AESL_inst_dft.temp_195_loc_channel_U.if_full_n;
    assign fifo_intf_196.fifo_rd_block = 0;
    assign fifo_intf_196.fifo_wr_block = 0;
    assign fifo_intf_196.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_196;
    csv_file_dump cstatus_csv_dumper_196;
    df_fifo_monitor fifo_monitor_196;
    df_fifo_intf fifo_intf_197(clock,reset);
    assign fifo_intf_197.rd_en = AESL_inst_dft.temp_196_loc_channel_U.if_read & AESL_inst_dft.temp_196_loc_channel_U.if_empty_n;
    assign fifo_intf_197.wr_en = AESL_inst_dft.temp_196_loc_channel_U.if_write & AESL_inst_dft.temp_196_loc_channel_U.if_full_n;
    assign fifo_intf_197.fifo_rd_block = 0;
    assign fifo_intf_197.fifo_wr_block = 0;
    assign fifo_intf_197.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_197;
    csv_file_dump cstatus_csv_dumper_197;
    df_fifo_monitor fifo_monitor_197;
    df_fifo_intf fifo_intf_198(clock,reset);
    assign fifo_intf_198.rd_en = AESL_inst_dft.temp_197_loc_channel_U.if_read & AESL_inst_dft.temp_197_loc_channel_U.if_empty_n;
    assign fifo_intf_198.wr_en = AESL_inst_dft.temp_197_loc_channel_U.if_write & AESL_inst_dft.temp_197_loc_channel_U.if_full_n;
    assign fifo_intf_198.fifo_rd_block = 0;
    assign fifo_intf_198.fifo_wr_block = 0;
    assign fifo_intf_198.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_198;
    csv_file_dump cstatus_csv_dumper_198;
    df_fifo_monitor fifo_monitor_198;
    df_fifo_intf fifo_intf_199(clock,reset);
    assign fifo_intf_199.rd_en = AESL_inst_dft.temp_198_loc_channel_U.if_read & AESL_inst_dft.temp_198_loc_channel_U.if_empty_n;
    assign fifo_intf_199.wr_en = AESL_inst_dft.temp_198_loc_channel_U.if_write & AESL_inst_dft.temp_198_loc_channel_U.if_full_n;
    assign fifo_intf_199.fifo_rd_block = 0;
    assign fifo_intf_199.fifo_wr_block = 0;
    assign fifo_intf_199.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_199;
    csv_file_dump cstatus_csv_dumper_199;
    df_fifo_monitor fifo_monitor_199;
    df_fifo_intf fifo_intf_200(clock,reset);
    assign fifo_intf_200.rd_en = AESL_inst_dft.temp_199_loc_channel_U.if_read & AESL_inst_dft.temp_199_loc_channel_U.if_empty_n;
    assign fifo_intf_200.wr_en = AESL_inst_dft.temp_199_loc_channel_U.if_write & AESL_inst_dft.temp_199_loc_channel_U.if_full_n;
    assign fifo_intf_200.fifo_rd_block = 0;
    assign fifo_intf_200.fifo_wr_block = 0;
    assign fifo_intf_200.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_200;
    csv_file_dump cstatus_csv_dumper_200;
    df_fifo_monitor fifo_monitor_200;
    df_fifo_intf fifo_intf_201(clock,reset);
    assign fifo_intf_201.rd_en = AESL_inst_dft.temp_200_loc_channel_U.if_read & AESL_inst_dft.temp_200_loc_channel_U.if_empty_n;
    assign fifo_intf_201.wr_en = AESL_inst_dft.temp_200_loc_channel_U.if_write & AESL_inst_dft.temp_200_loc_channel_U.if_full_n;
    assign fifo_intf_201.fifo_rd_block = 0;
    assign fifo_intf_201.fifo_wr_block = 0;
    assign fifo_intf_201.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_201;
    csv_file_dump cstatus_csv_dumper_201;
    df_fifo_monitor fifo_monitor_201;
    df_fifo_intf fifo_intf_202(clock,reset);
    assign fifo_intf_202.rd_en = AESL_inst_dft.temp_201_loc_channel_U.if_read & AESL_inst_dft.temp_201_loc_channel_U.if_empty_n;
    assign fifo_intf_202.wr_en = AESL_inst_dft.temp_201_loc_channel_U.if_write & AESL_inst_dft.temp_201_loc_channel_U.if_full_n;
    assign fifo_intf_202.fifo_rd_block = 0;
    assign fifo_intf_202.fifo_wr_block = 0;
    assign fifo_intf_202.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_202;
    csv_file_dump cstatus_csv_dumper_202;
    df_fifo_monitor fifo_monitor_202;
    df_fifo_intf fifo_intf_203(clock,reset);
    assign fifo_intf_203.rd_en = AESL_inst_dft.temp_202_loc_channel_U.if_read & AESL_inst_dft.temp_202_loc_channel_U.if_empty_n;
    assign fifo_intf_203.wr_en = AESL_inst_dft.temp_202_loc_channel_U.if_write & AESL_inst_dft.temp_202_loc_channel_U.if_full_n;
    assign fifo_intf_203.fifo_rd_block = 0;
    assign fifo_intf_203.fifo_wr_block = 0;
    assign fifo_intf_203.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_203;
    csv_file_dump cstatus_csv_dumper_203;
    df_fifo_monitor fifo_monitor_203;
    df_fifo_intf fifo_intf_204(clock,reset);
    assign fifo_intf_204.rd_en = AESL_inst_dft.temp_203_loc_channel_U.if_read & AESL_inst_dft.temp_203_loc_channel_U.if_empty_n;
    assign fifo_intf_204.wr_en = AESL_inst_dft.temp_203_loc_channel_U.if_write & AESL_inst_dft.temp_203_loc_channel_U.if_full_n;
    assign fifo_intf_204.fifo_rd_block = 0;
    assign fifo_intf_204.fifo_wr_block = 0;
    assign fifo_intf_204.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_204;
    csv_file_dump cstatus_csv_dumper_204;
    df_fifo_monitor fifo_monitor_204;
    df_fifo_intf fifo_intf_205(clock,reset);
    assign fifo_intf_205.rd_en = AESL_inst_dft.temp_204_loc_channel_U.if_read & AESL_inst_dft.temp_204_loc_channel_U.if_empty_n;
    assign fifo_intf_205.wr_en = AESL_inst_dft.temp_204_loc_channel_U.if_write & AESL_inst_dft.temp_204_loc_channel_U.if_full_n;
    assign fifo_intf_205.fifo_rd_block = 0;
    assign fifo_intf_205.fifo_wr_block = 0;
    assign fifo_intf_205.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_205;
    csv_file_dump cstatus_csv_dumper_205;
    df_fifo_monitor fifo_monitor_205;
    df_fifo_intf fifo_intf_206(clock,reset);
    assign fifo_intf_206.rd_en = AESL_inst_dft.temp_205_loc_channel_U.if_read & AESL_inst_dft.temp_205_loc_channel_U.if_empty_n;
    assign fifo_intf_206.wr_en = AESL_inst_dft.temp_205_loc_channel_U.if_write & AESL_inst_dft.temp_205_loc_channel_U.if_full_n;
    assign fifo_intf_206.fifo_rd_block = 0;
    assign fifo_intf_206.fifo_wr_block = 0;
    assign fifo_intf_206.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_206;
    csv_file_dump cstatus_csv_dumper_206;
    df_fifo_monitor fifo_monitor_206;
    df_fifo_intf fifo_intf_207(clock,reset);
    assign fifo_intf_207.rd_en = AESL_inst_dft.temp_206_loc_channel_U.if_read & AESL_inst_dft.temp_206_loc_channel_U.if_empty_n;
    assign fifo_intf_207.wr_en = AESL_inst_dft.temp_206_loc_channel_U.if_write & AESL_inst_dft.temp_206_loc_channel_U.if_full_n;
    assign fifo_intf_207.fifo_rd_block = 0;
    assign fifo_intf_207.fifo_wr_block = 0;
    assign fifo_intf_207.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_207;
    csv_file_dump cstatus_csv_dumper_207;
    df_fifo_monitor fifo_monitor_207;
    df_fifo_intf fifo_intf_208(clock,reset);
    assign fifo_intf_208.rd_en = AESL_inst_dft.temp_207_loc_channel_U.if_read & AESL_inst_dft.temp_207_loc_channel_U.if_empty_n;
    assign fifo_intf_208.wr_en = AESL_inst_dft.temp_207_loc_channel_U.if_write & AESL_inst_dft.temp_207_loc_channel_U.if_full_n;
    assign fifo_intf_208.fifo_rd_block = 0;
    assign fifo_intf_208.fifo_wr_block = 0;
    assign fifo_intf_208.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_208;
    csv_file_dump cstatus_csv_dumper_208;
    df_fifo_monitor fifo_monitor_208;
    df_fifo_intf fifo_intf_209(clock,reset);
    assign fifo_intf_209.rd_en = AESL_inst_dft.temp_208_loc_channel_U.if_read & AESL_inst_dft.temp_208_loc_channel_U.if_empty_n;
    assign fifo_intf_209.wr_en = AESL_inst_dft.temp_208_loc_channel_U.if_write & AESL_inst_dft.temp_208_loc_channel_U.if_full_n;
    assign fifo_intf_209.fifo_rd_block = 0;
    assign fifo_intf_209.fifo_wr_block = 0;
    assign fifo_intf_209.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_209;
    csv_file_dump cstatus_csv_dumper_209;
    df_fifo_monitor fifo_monitor_209;
    df_fifo_intf fifo_intf_210(clock,reset);
    assign fifo_intf_210.rd_en = AESL_inst_dft.temp_209_loc_channel_U.if_read & AESL_inst_dft.temp_209_loc_channel_U.if_empty_n;
    assign fifo_intf_210.wr_en = AESL_inst_dft.temp_209_loc_channel_U.if_write & AESL_inst_dft.temp_209_loc_channel_U.if_full_n;
    assign fifo_intf_210.fifo_rd_block = 0;
    assign fifo_intf_210.fifo_wr_block = 0;
    assign fifo_intf_210.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_210;
    csv_file_dump cstatus_csv_dumper_210;
    df_fifo_monitor fifo_monitor_210;
    df_fifo_intf fifo_intf_211(clock,reset);
    assign fifo_intf_211.rd_en = AESL_inst_dft.temp_210_loc_channel_U.if_read & AESL_inst_dft.temp_210_loc_channel_U.if_empty_n;
    assign fifo_intf_211.wr_en = AESL_inst_dft.temp_210_loc_channel_U.if_write & AESL_inst_dft.temp_210_loc_channel_U.if_full_n;
    assign fifo_intf_211.fifo_rd_block = 0;
    assign fifo_intf_211.fifo_wr_block = 0;
    assign fifo_intf_211.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_211;
    csv_file_dump cstatus_csv_dumper_211;
    df_fifo_monitor fifo_monitor_211;
    df_fifo_intf fifo_intf_212(clock,reset);
    assign fifo_intf_212.rd_en = AESL_inst_dft.temp_211_loc_channel_U.if_read & AESL_inst_dft.temp_211_loc_channel_U.if_empty_n;
    assign fifo_intf_212.wr_en = AESL_inst_dft.temp_211_loc_channel_U.if_write & AESL_inst_dft.temp_211_loc_channel_U.if_full_n;
    assign fifo_intf_212.fifo_rd_block = 0;
    assign fifo_intf_212.fifo_wr_block = 0;
    assign fifo_intf_212.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_212;
    csv_file_dump cstatus_csv_dumper_212;
    df_fifo_monitor fifo_monitor_212;
    df_fifo_intf fifo_intf_213(clock,reset);
    assign fifo_intf_213.rd_en = AESL_inst_dft.temp_212_loc_channel_U.if_read & AESL_inst_dft.temp_212_loc_channel_U.if_empty_n;
    assign fifo_intf_213.wr_en = AESL_inst_dft.temp_212_loc_channel_U.if_write & AESL_inst_dft.temp_212_loc_channel_U.if_full_n;
    assign fifo_intf_213.fifo_rd_block = 0;
    assign fifo_intf_213.fifo_wr_block = 0;
    assign fifo_intf_213.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_213;
    csv_file_dump cstatus_csv_dumper_213;
    df_fifo_monitor fifo_monitor_213;
    df_fifo_intf fifo_intf_214(clock,reset);
    assign fifo_intf_214.rd_en = AESL_inst_dft.temp_213_loc_channel_U.if_read & AESL_inst_dft.temp_213_loc_channel_U.if_empty_n;
    assign fifo_intf_214.wr_en = AESL_inst_dft.temp_213_loc_channel_U.if_write & AESL_inst_dft.temp_213_loc_channel_U.if_full_n;
    assign fifo_intf_214.fifo_rd_block = 0;
    assign fifo_intf_214.fifo_wr_block = 0;
    assign fifo_intf_214.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_214;
    csv_file_dump cstatus_csv_dumper_214;
    df_fifo_monitor fifo_monitor_214;
    df_fifo_intf fifo_intf_215(clock,reset);
    assign fifo_intf_215.rd_en = AESL_inst_dft.temp_214_loc_channel_U.if_read & AESL_inst_dft.temp_214_loc_channel_U.if_empty_n;
    assign fifo_intf_215.wr_en = AESL_inst_dft.temp_214_loc_channel_U.if_write & AESL_inst_dft.temp_214_loc_channel_U.if_full_n;
    assign fifo_intf_215.fifo_rd_block = 0;
    assign fifo_intf_215.fifo_wr_block = 0;
    assign fifo_intf_215.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_215;
    csv_file_dump cstatus_csv_dumper_215;
    df_fifo_monitor fifo_monitor_215;
    df_fifo_intf fifo_intf_216(clock,reset);
    assign fifo_intf_216.rd_en = AESL_inst_dft.temp_215_loc_channel_U.if_read & AESL_inst_dft.temp_215_loc_channel_U.if_empty_n;
    assign fifo_intf_216.wr_en = AESL_inst_dft.temp_215_loc_channel_U.if_write & AESL_inst_dft.temp_215_loc_channel_U.if_full_n;
    assign fifo_intf_216.fifo_rd_block = 0;
    assign fifo_intf_216.fifo_wr_block = 0;
    assign fifo_intf_216.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_216;
    csv_file_dump cstatus_csv_dumper_216;
    df_fifo_monitor fifo_monitor_216;
    df_fifo_intf fifo_intf_217(clock,reset);
    assign fifo_intf_217.rd_en = AESL_inst_dft.temp_216_loc_channel_U.if_read & AESL_inst_dft.temp_216_loc_channel_U.if_empty_n;
    assign fifo_intf_217.wr_en = AESL_inst_dft.temp_216_loc_channel_U.if_write & AESL_inst_dft.temp_216_loc_channel_U.if_full_n;
    assign fifo_intf_217.fifo_rd_block = 0;
    assign fifo_intf_217.fifo_wr_block = 0;
    assign fifo_intf_217.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_217;
    csv_file_dump cstatus_csv_dumper_217;
    df_fifo_monitor fifo_monitor_217;
    df_fifo_intf fifo_intf_218(clock,reset);
    assign fifo_intf_218.rd_en = AESL_inst_dft.temp_217_loc_channel_U.if_read & AESL_inst_dft.temp_217_loc_channel_U.if_empty_n;
    assign fifo_intf_218.wr_en = AESL_inst_dft.temp_217_loc_channel_U.if_write & AESL_inst_dft.temp_217_loc_channel_U.if_full_n;
    assign fifo_intf_218.fifo_rd_block = 0;
    assign fifo_intf_218.fifo_wr_block = 0;
    assign fifo_intf_218.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_218;
    csv_file_dump cstatus_csv_dumper_218;
    df_fifo_monitor fifo_monitor_218;
    df_fifo_intf fifo_intf_219(clock,reset);
    assign fifo_intf_219.rd_en = AESL_inst_dft.temp_218_loc_channel_U.if_read & AESL_inst_dft.temp_218_loc_channel_U.if_empty_n;
    assign fifo_intf_219.wr_en = AESL_inst_dft.temp_218_loc_channel_U.if_write & AESL_inst_dft.temp_218_loc_channel_U.if_full_n;
    assign fifo_intf_219.fifo_rd_block = 0;
    assign fifo_intf_219.fifo_wr_block = 0;
    assign fifo_intf_219.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_219;
    csv_file_dump cstatus_csv_dumper_219;
    df_fifo_monitor fifo_monitor_219;
    df_fifo_intf fifo_intf_220(clock,reset);
    assign fifo_intf_220.rd_en = AESL_inst_dft.temp_219_loc_channel_U.if_read & AESL_inst_dft.temp_219_loc_channel_U.if_empty_n;
    assign fifo_intf_220.wr_en = AESL_inst_dft.temp_219_loc_channel_U.if_write & AESL_inst_dft.temp_219_loc_channel_U.if_full_n;
    assign fifo_intf_220.fifo_rd_block = 0;
    assign fifo_intf_220.fifo_wr_block = 0;
    assign fifo_intf_220.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_220;
    csv_file_dump cstatus_csv_dumper_220;
    df_fifo_monitor fifo_monitor_220;
    df_fifo_intf fifo_intf_221(clock,reset);
    assign fifo_intf_221.rd_en = AESL_inst_dft.temp_220_loc_channel_U.if_read & AESL_inst_dft.temp_220_loc_channel_U.if_empty_n;
    assign fifo_intf_221.wr_en = AESL_inst_dft.temp_220_loc_channel_U.if_write & AESL_inst_dft.temp_220_loc_channel_U.if_full_n;
    assign fifo_intf_221.fifo_rd_block = 0;
    assign fifo_intf_221.fifo_wr_block = 0;
    assign fifo_intf_221.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_221;
    csv_file_dump cstatus_csv_dumper_221;
    df_fifo_monitor fifo_monitor_221;
    df_fifo_intf fifo_intf_222(clock,reset);
    assign fifo_intf_222.rd_en = AESL_inst_dft.temp_221_loc_channel_U.if_read & AESL_inst_dft.temp_221_loc_channel_U.if_empty_n;
    assign fifo_intf_222.wr_en = AESL_inst_dft.temp_221_loc_channel_U.if_write & AESL_inst_dft.temp_221_loc_channel_U.if_full_n;
    assign fifo_intf_222.fifo_rd_block = 0;
    assign fifo_intf_222.fifo_wr_block = 0;
    assign fifo_intf_222.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_222;
    csv_file_dump cstatus_csv_dumper_222;
    df_fifo_monitor fifo_monitor_222;
    df_fifo_intf fifo_intf_223(clock,reset);
    assign fifo_intf_223.rd_en = AESL_inst_dft.temp_222_loc_channel_U.if_read & AESL_inst_dft.temp_222_loc_channel_U.if_empty_n;
    assign fifo_intf_223.wr_en = AESL_inst_dft.temp_222_loc_channel_U.if_write & AESL_inst_dft.temp_222_loc_channel_U.if_full_n;
    assign fifo_intf_223.fifo_rd_block = 0;
    assign fifo_intf_223.fifo_wr_block = 0;
    assign fifo_intf_223.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_223;
    csv_file_dump cstatus_csv_dumper_223;
    df_fifo_monitor fifo_monitor_223;
    df_fifo_intf fifo_intf_224(clock,reset);
    assign fifo_intf_224.rd_en = AESL_inst_dft.temp_223_loc_channel_U.if_read & AESL_inst_dft.temp_223_loc_channel_U.if_empty_n;
    assign fifo_intf_224.wr_en = AESL_inst_dft.temp_223_loc_channel_U.if_write & AESL_inst_dft.temp_223_loc_channel_U.if_full_n;
    assign fifo_intf_224.fifo_rd_block = 0;
    assign fifo_intf_224.fifo_wr_block = 0;
    assign fifo_intf_224.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_224;
    csv_file_dump cstatus_csv_dumper_224;
    df_fifo_monitor fifo_monitor_224;
    df_fifo_intf fifo_intf_225(clock,reset);
    assign fifo_intf_225.rd_en = AESL_inst_dft.temp_224_loc_channel_U.if_read & AESL_inst_dft.temp_224_loc_channel_U.if_empty_n;
    assign fifo_intf_225.wr_en = AESL_inst_dft.temp_224_loc_channel_U.if_write & AESL_inst_dft.temp_224_loc_channel_U.if_full_n;
    assign fifo_intf_225.fifo_rd_block = 0;
    assign fifo_intf_225.fifo_wr_block = 0;
    assign fifo_intf_225.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_225;
    csv_file_dump cstatus_csv_dumper_225;
    df_fifo_monitor fifo_monitor_225;
    df_fifo_intf fifo_intf_226(clock,reset);
    assign fifo_intf_226.rd_en = AESL_inst_dft.temp_225_loc_channel_U.if_read & AESL_inst_dft.temp_225_loc_channel_U.if_empty_n;
    assign fifo_intf_226.wr_en = AESL_inst_dft.temp_225_loc_channel_U.if_write & AESL_inst_dft.temp_225_loc_channel_U.if_full_n;
    assign fifo_intf_226.fifo_rd_block = 0;
    assign fifo_intf_226.fifo_wr_block = 0;
    assign fifo_intf_226.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_226;
    csv_file_dump cstatus_csv_dumper_226;
    df_fifo_monitor fifo_monitor_226;
    df_fifo_intf fifo_intf_227(clock,reset);
    assign fifo_intf_227.rd_en = AESL_inst_dft.temp_226_loc_channel_U.if_read & AESL_inst_dft.temp_226_loc_channel_U.if_empty_n;
    assign fifo_intf_227.wr_en = AESL_inst_dft.temp_226_loc_channel_U.if_write & AESL_inst_dft.temp_226_loc_channel_U.if_full_n;
    assign fifo_intf_227.fifo_rd_block = 0;
    assign fifo_intf_227.fifo_wr_block = 0;
    assign fifo_intf_227.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_227;
    csv_file_dump cstatus_csv_dumper_227;
    df_fifo_monitor fifo_monitor_227;
    df_fifo_intf fifo_intf_228(clock,reset);
    assign fifo_intf_228.rd_en = AESL_inst_dft.temp_227_loc_channel_U.if_read & AESL_inst_dft.temp_227_loc_channel_U.if_empty_n;
    assign fifo_intf_228.wr_en = AESL_inst_dft.temp_227_loc_channel_U.if_write & AESL_inst_dft.temp_227_loc_channel_U.if_full_n;
    assign fifo_intf_228.fifo_rd_block = 0;
    assign fifo_intf_228.fifo_wr_block = 0;
    assign fifo_intf_228.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_228;
    csv_file_dump cstatus_csv_dumper_228;
    df_fifo_monitor fifo_monitor_228;
    df_fifo_intf fifo_intf_229(clock,reset);
    assign fifo_intf_229.rd_en = AESL_inst_dft.temp_228_loc_channel_U.if_read & AESL_inst_dft.temp_228_loc_channel_U.if_empty_n;
    assign fifo_intf_229.wr_en = AESL_inst_dft.temp_228_loc_channel_U.if_write & AESL_inst_dft.temp_228_loc_channel_U.if_full_n;
    assign fifo_intf_229.fifo_rd_block = 0;
    assign fifo_intf_229.fifo_wr_block = 0;
    assign fifo_intf_229.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_229;
    csv_file_dump cstatus_csv_dumper_229;
    df_fifo_monitor fifo_monitor_229;
    df_fifo_intf fifo_intf_230(clock,reset);
    assign fifo_intf_230.rd_en = AESL_inst_dft.temp_229_loc_channel_U.if_read & AESL_inst_dft.temp_229_loc_channel_U.if_empty_n;
    assign fifo_intf_230.wr_en = AESL_inst_dft.temp_229_loc_channel_U.if_write & AESL_inst_dft.temp_229_loc_channel_U.if_full_n;
    assign fifo_intf_230.fifo_rd_block = 0;
    assign fifo_intf_230.fifo_wr_block = 0;
    assign fifo_intf_230.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_230;
    csv_file_dump cstatus_csv_dumper_230;
    df_fifo_monitor fifo_monitor_230;
    df_fifo_intf fifo_intf_231(clock,reset);
    assign fifo_intf_231.rd_en = AESL_inst_dft.temp_230_loc_channel_U.if_read & AESL_inst_dft.temp_230_loc_channel_U.if_empty_n;
    assign fifo_intf_231.wr_en = AESL_inst_dft.temp_230_loc_channel_U.if_write & AESL_inst_dft.temp_230_loc_channel_U.if_full_n;
    assign fifo_intf_231.fifo_rd_block = 0;
    assign fifo_intf_231.fifo_wr_block = 0;
    assign fifo_intf_231.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_231;
    csv_file_dump cstatus_csv_dumper_231;
    df_fifo_monitor fifo_monitor_231;
    df_fifo_intf fifo_intf_232(clock,reset);
    assign fifo_intf_232.rd_en = AESL_inst_dft.temp_231_loc_channel_U.if_read & AESL_inst_dft.temp_231_loc_channel_U.if_empty_n;
    assign fifo_intf_232.wr_en = AESL_inst_dft.temp_231_loc_channel_U.if_write & AESL_inst_dft.temp_231_loc_channel_U.if_full_n;
    assign fifo_intf_232.fifo_rd_block = 0;
    assign fifo_intf_232.fifo_wr_block = 0;
    assign fifo_intf_232.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_232;
    csv_file_dump cstatus_csv_dumper_232;
    df_fifo_monitor fifo_monitor_232;
    df_fifo_intf fifo_intf_233(clock,reset);
    assign fifo_intf_233.rd_en = AESL_inst_dft.temp_232_loc_channel_U.if_read & AESL_inst_dft.temp_232_loc_channel_U.if_empty_n;
    assign fifo_intf_233.wr_en = AESL_inst_dft.temp_232_loc_channel_U.if_write & AESL_inst_dft.temp_232_loc_channel_U.if_full_n;
    assign fifo_intf_233.fifo_rd_block = 0;
    assign fifo_intf_233.fifo_wr_block = 0;
    assign fifo_intf_233.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_233;
    csv_file_dump cstatus_csv_dumper_233;
    df_fifo_monitor fifo_monitor_233;
    df_fifo_intf fifo_intf_234(clock,reset);
    assign fifo_intf_234.rd_en = AESL_inst_dft.temp_233_loc_channel_U.if_read & AESL_inst_dft.temp_233_loc_channel_U.if_empty_n;
    assign fifo_intf_234.wr_en = AESL_inst_dft.temp_233_loc_channel_U.if_write & AESL_inst_dft.temp_233_loc_channel_U.if_full_n;
    assign fifo_intf_234.fifo_rd_block = 0;
    assign fifo_intf_234.fifo_wr_block = 0;
    assign fifo_intf_234.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_234;
    csv_file_dump cstatus_csv_dumper_234;
    df_fifo_monitor fifo_monitor_234;
    df_fifo_intf fifo_intf_235(clock,reset);
    assign fifo_intf_235.rd_en = AESL_inst_dft.temp_234_loc_channel_U.if_read & AESL_inst_dft.temp_234_loc_channel_U.if_empty_n;
    assign fifo_intf_235.wr_en = AESL_inst_dft.temp_234_loc_channel_U.if_write & AESL_inst_dft.temp_234_loc_channel_U.if_full_n;
    assign fifo_intf_235.fifo_rd_block = 0;
    assign fifo_intf_235.fifo_wr_block = 0;
    assign fifo_intf_235.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_235;
    csv_file_dump cstatus_csv_dumper_235;
    df_fifo_monitor fifo_monitor_235;
    df_fifo_intf fifo_intf_236(clock,reset);
    assign fifo_intf_236.rd_en = AESL_inst_dft.temp_235_loc_channel_U.if_read & AESL_inst_dft.temp_235_loc_channel_U.if_empty_n;
    assign fifo_intf_236.wr_en = AESL_inst_dft.temp_235_loc_channel_U.if_write & AESL_inst_dft.temp_235_loc_channel_U.if_full_n;
    assign fifo_intf_236.fifo_rd_block = 0;
    assign fifo_intf_236.fifo_wr_block = 0;
    assign fifo_intf_236.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_236;
    csv_file_dump cstatus_csv_dumper_236;
    df_fifo_monitor fifo_monitor_236;
    df_fifo_intf fifo_intf_237(clock,reset);
    assign fifo_intf_237.rd_en = AESL_inst_dft.temp_236_loc_channel_U.if_read & AESL_inst_dft.temp_236_loc_channel_U.if_empty_n;
    assign fifo_intf_237.wr_en = AESL_inst_dft.temp_236_loc_channel_U.if_write & AESL_inst_dft.temp_236_loc_channel_U.if_full_n;
    assign fifo_intf_237.fifo_rd_block = 0;
    assign fifo_intf_237.fifo_wr_block = 0;
    assign fifo_intf_237.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_237;
    csv_file_dump cstatus_csv_dumper_237;
    df_fifo_monitor fifo_monitor_237;
    df_fifo_intf fifo_intf_238(clock,reset);
    assign fifo_intf_238.rd_en = AESL_inst_dft.temp_237_loc_channel_U.if_read & AESL_inst_dft.temp_237_loc_channel_U.if_empty_n;
    assign fifo_intf_238.wr_en = AESL_inst_dft.temp_237_loc_channel_U.if_write & AESL_inst_dft.temp_237_loc_channel_U.if_full_n;
    assign fifo_intf_238.fifo_rd_block = 0;
    assign fifo_intf_238.fifo_wr_block = 0;
    assign fifo_intf_238.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_238;
    csv_file_dump cstatus_csv_dumper_238;
    df_fifo_monitor fifo_monitor_238;
    df_fifo_intf fifo_intf_239(clock,reset);
    assign fifo_intf_239.rd_en = AESL_inst_dft.temp_238_loc_channel_U.if_read & AESL_inst_dft.temp_238_loc_channel_U.if_empty_n;
    assign fifo_intf_239.wr_en = AESL_inst_dft.temp_238_loc_channel_U.if_write & AESL_inst_dft.temp_238_loc_channel_U.if_full_n;
    assign fifo_intf_239.fifo_rd_block = 0;
    assign fifo_intf_239.fifo_wr_block = 0;
    assign fifo_intf_239.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_239;
    csv_file_dump cstatus_csv_dumper_239;
    df_fifo_monitor fifo_monitor_239;
    df_fifo_intf fifo_intf_240(clock,reset);
    assign fifo_intf_240.rd_en = AESL_inst_dft.temp_239_loc_channel_U.if_read & AESL_inst_dft.temp_239_loc_channel_U.if_empty_n;
    assign fifo_intf_240.wr_en = AESL_inst_dft.temp_239_loc_channel_U.if_write & AESL_inst_dft.temp_239_loc_channel_U.if_full_n;
    assign fifo_intf_240.fifo_rd_block = 0;
    assign fifo_intf_240.fifo_wr_block = 0;
    assign fifo_intf_240.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_240;
    csv_file_dump cstatus_csv_dumper_240;
    df_fifo_monitor fifo_monitor_240;
    df_fifo_intf fifo_intf_241(clock,reset);
    assign fifo_intf_241.rd_en = AESL_inst_dft.temp_240_loc_channel_U.if_read & AESL_inst_dft.temp_240_loc_channel_U.if_empty_n;
    assign fifo_intf_241.wr_en = AESL_inst_dft.temp_240_loc_channel_U.if_write & AESL_inst_dft.temp_240_loc_channel_U.if_full_n;
    assign fifo_intf_241.fifo_rd_block = 0;
    assign fifo_intf_241.fifo_wr_block = 0;
    assign fifo_intf_241.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_241;
    csv_file_dump cstatus_csv_dumper_241;
    df_fifo_monitor fifo_monitor_241;
    df_fifo_intf fifo_intf_242(clock,reset);
    assign fifo_intf_242.rd_en = AESL_inst_dft.temp_241_loc_channel_U.if_read & AESL_inst_dft.temp_241_loc_channel_U.if_empty_n;
    assign fifo_intf_242.wr_en = AESL_inst_dft.temp_241_loc_channel_U.if_write & AESL_inst_dft.temp_241_loc_channel_U.if_full_n;
    assign fifo_intf_242.fifo_rd_block = 0;
    assign fifo_intf_242.fifo_wr_block = 0;
    assign fifo_intf_242.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_242;
    csv_file_dump cstatus_csv_dumper_242;
    df_fifo_monitor fifo_monitor_242;
    df_fifo_intf fifo_intf_243(clock,reset);
    assign fifo_intf_243.rd_en = AESL_inst_dft.temp_242_loc_channel_U.if_read & AESL_inst_dft.temp_242_loc_channel_U.if_empty_n;
    assign fifo_intf_243.wr_en = AESL_inst_dft.temp_242_loc_channel_U.if_write & AESL_inst_dft.temp_242_loc_channel_U.if_full_n;
    assign fifo_intf_243.fifo_rd_block = 0;
    assign fifo_intf_243.fifo_wr_block = 0;
    assign fifo_intf_243.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_243;
    csv_file_dump cstatus_csv_dumper_243;
    df_fifo_monitor fifo_monitor_243;
    df_fifo_intf fifo_intf_244(clock,reset);
    assign fifo_intf_244.rd_en = AESL_inst_dft.temp_243_loc_channel_U.if_read & AESL_inst_dft.temp_243_loc_channel_U.if_empty_n;
    assign fifo_intf_244.wr_en = AESL_inst_dft.temp_243_loc_channel_U.if_write & AESL_inst_dft.temp_243_loc_channel_U.if_full_n;
    assign fifo_intf_244.fifo_rd_block = 0;
    assign fifo_intf_244.fifo_wr_block = 0;
    assign fifo_intf_244.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_244;
    csv_file_dump cstatus_csv_dumper_244;
    df_fifo_monitor fifo_monitor_244;
    df_fifo_intf fifo_intf_245(clock,reset);
    assign fifo_intf_245.rd_en = AESL_inst_dft.temp_244_loc_channel_U.if_read & AESL_inst_dft.temp_244_loc_channel_U.if_empty_n;
    assign fifo_intf_245.wr_en = AESL_inst_dft.temp_244_loc_channel_U.if_write & AESL_inst_dft.temp_244_loc_channel_U.if_full_n;
    assign fifo_intf_245.fifo_rd_block = 0;
    assign fifo_intf_245.fifo_wr_block = 0;
    assign fifo_intf_245.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_245;
    csv_file_dump cstatus_csv_dumper_245;
    df_fifo_monitor fifo_monitor_245;
    df_fifo_intf fifo_intf_246(clock,reset);
    assign fifo_intf_246.rd_en = AESL_inst_dft.temp_245_loc_channel_U.if_read & AESL_inst_dft.temp_245_loc_channel_U.if_empty_n;
    assign fifo_intf_246.wr_en = AESL_inst_dft.temp_245_loc_channel_U.if_write & AESL_inst_dft.temp_245_loc_channel_U.if_full_n;
    assign fifo_intf_246.fifo_rd_block = 0;
    assign fifo_intf_246.fifo_wr_block = 0;
    assign fifo_intf_246.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_246;
    csv_file_dump cstatus_csv_dumper_246;
    df_fifo_monitor fifo_monitor_246;
    df_fifo_intf fifo_intf_247(clock,reset);
    assign fifo_intf_247.rd_en = AESL_inst_dft.temp_246_loc_channel_U.if_read & AESL_inst_dft.temp_246_loc_channel_U.if_empty_n;
    assign fifo_intf_247.wr_en = AESL_inst_dft.temp_246_loc_channel_U.if_write & AESL_inst_dft.temp_246_loc_channel_U.if_full_n;
    assign fifo_intf_247.fifo_rd_block = 0;
    assign fifo_intf_247.fifo_wr_block = 0;
    assign fifo_intf_247.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_247;
    csv_file_dump cstatus_csv_dumper_247;
    df_fifo_monitor fifo_monitor_247;
    df_fifo_intf fifo_intf_248(clock,reset);
    assign fifo_intf_248.rd_en = AESL_inst_dft.temp_247_loc_channel_U.if_read & AESL_inst_dft.temp_247_loc_channel_U.if_empty_n;
    assign fifo_intf_248.wr_en = AESL_inst_dft.temp_247_loc_channel_U.if_write & AESL_inst_dft.temp_247_loc_channel_U.if_full_n;
    assign fifo_intf_248.fifo_rd_block = 0;
    assign fifo_intf_248.fifo_wr_block = 0;
    assign fifo_intf_248.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_248;
    csv_file_dump cstatus_csv_dumper_248;
    df_fifo_monitor fifo_monitor_248;
    df_fifo_intf fifo_intf_249(clock,reset);
    assign fifo_intf_249.rd_en = AESL_inst_dft.temp_248_loc_channel_U.if_read & AESL_inst_dft.temp_248_loc_channel_U.if_empty_n;
    assign fifo_intf_249.wr_en = AESL_inst_dft.temp_248_loc_channel_U.if_write & AESL_inst_dft.temp_248_loc_channel_U.if_full_n;
    assign fifo_intf_249.fifo_rd_block = 0;
    assign fifo_intf_249.fifo_wr_block = 0;
    assign fifo_intf_249.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_249;
    csv_file_dump cstatus_csv_dumper_249;
    df_fifo_monitor fifo_monitor_249;
    df_fifo_intf fifo_intf_250(clock,reset);
    assign fifo_intf_250.rd_en = AESL_inst_dft.temp_249_loc_channel_U.if_read & AESL_inst_dft.temp_249_loc_channel_U.if_empty_n;
    assign fifo_intf_250.wr_en = AESL_inst_dft.temp_249_loc_channel_U.if_write & AESL_inst_dft.temp_249_loc_channel_U.if_full_n;
    assign fifo_intf_250.fifo_rd_block = 0;
    assign fifo_intf_250.fifo_wr_block = 0;
    assign fifo_intf_250.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_250;
    csv_file_dump cstatus_csv_dumper_250;
    df_fifo_monitor fifo_monitor_250;
    df_fifo_intf fifo_intf_251(clock,reset);
    assign fifo_intf_251.rd_en = AESL_inst_dft.temp_250_loc_channel_U.if_read & AESL_inst_dft.temp_250_loc_channel_U.if_empty_n;
    assign fifo_intf_251.wr_en = AESL_inst_dft.temp_250_loc_channel_U.if_write & AESL_inst_dft.temp_250_loc_channel_U.if_full_n;
    assign fifo_intf_251.fifo_rd_block = 0;
    assign fifo_intf_251.fifo_wr_block = 0;
    assign fifo_intf_251.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_251;
    csv_file_dump cstatus_csv_dumper_251;
    df_fifo_monitor fifo_monitor_251;
    df_fifo_intf fifo_intf_252(clock,reset);
    assign fifo_intf_252.rd_en = AESL_inst_dft.temp_251_loc_channel_U.if_read & AESL_inst_dft.temp_251_loc_channel_U.if_empty_n;
    assign fifo_intf_252.wr_en = AESL_inst_dft.temp_251_loc_channel_U.if_write & AESL_inst_dft.temp_251_loc_channel_U.if_full_n;
    assign fifo_intf_252.fifo_rd_block = 0;
    assign fifo_intf_252.fifo_wr_block = 0;
    assign fifo_intf_252.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_252;
    csv_file_dump cstatus_csv_dumper_252;
    df_fifo_monitor fifo_monitor_252;
    df_fifo_intf fifo_intf_253(clock,reset);
    assign fifo_intf_253.rd_en = AESL_inst_dft.temp_252_loc_channel_U.if_read & AESL_inst_dft.temp_252_loc_channel_U.if_empty_n;
    assign fifo_intf_253.wr_en = AESL_inst_dft.temp_252_loc_channel_U.if_write & AESL_inst_dft.temp_252_loc_channel_U.if_full_n;
    assign fifo_intf_253.fifo_rd_block = 0;
    assign fifo_intf_253.fifo_wr_block = 0;
    assign fifo_intf_253.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_253;
    csv_file_dump cstatus_csv_dumper_253;
    df_fifo_monitor fifo_monitor_253;
    df_fifo_intf fifo_intf_254(clock,reset);
    assign fifo_intf_254.rd_en = AESL_inst_dft.temp_253_loc_channel_U.if_read & AESL_inst_dft.temp_253_loc_channel_U.if_empty_n;
    assign fifo_intf_254.wr_en = AESL_inst_dft.temp_253_loc_channel_U.if_write & AESL_inst_dft.temp_253_loc_channel_U.if_full_n;
    assign fifo_intf_254.fifo_rd_block = 0;
    assign fifo_intf_254.fifo_wr_block = 0;
    assign fifo_intf_254.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_254;
    csv_file_dump cstatus_csv_dumper_254;
    df_fifo_monitor fifo_monitor_254;
    df_fifo_intf fifo_intf_255(clock,reset);
    assign fifo_intf_255.rd_en = AESL_inst_dft.temp_254_loc_channel_U.if_read & AESL_inst_dft.temp_254_loc_channel_U.if_empty_n;
    assign fifo_intf_255.wr_en = AESL_inst_dft.temp_254_loc_channel_U.if_write & AESL_inst_dft.temp_254_loc_channel_U.if_full_n;
    assign fifo_intf_255.fifo_rd_block = 0;
    assign fifo_intf_255.fifo_wr_block = 0;
    assign fifo_intf_255.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_255;
    csv_file_dump cstatus_csv_dumper_255;
    df_fifo_monitor fifo_monitor_255;
    df_fifo_intf fifo_intf_256(clock,reset);
    assign fifo_intf_256.rd_en = AESL_inst_dft.temp_255_loc_channel_U.if_read & AESL_inst_dft.temp_255_loc_channel_U.if_empty_n;
    assign fifo_intf_256.wr_en = AESL_inst_dft.temp_255_loc_channel_U.if_write & AESL_inst_dft.temp_255_loc_channel_U.if_full_n;
    assign fifo_intf_256.fifo_rd_block = 0;
    assign fifo_intf_256.fifo_wr_block = 0;
    assign fifo_intf_256.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_256;
    csv_file_dump cstatus_csv_dumper_256;
    df_fifo_monitor fifo_monitor_256;

logic region_0_idle;
logic [31:0] region_0_start_cnt;
logic [31:0] region_0_done_cnt;
assign region_0_idle = (region_0_start_cnt == region_0_done_cnt) && AESL_inst_dft.ap_start == 1'b0 ;
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_start_cnt <= 32'h0;
    else if (AESL_inst_dft.ap_start == 1'b1 && AESL_inst_dft.ap_ready == 1'b1)
        region_0_start_cnt <= region_0_start_cnt + 32'h1;
    else;
end
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_done_cnt <= 32'h0;
    else if (AESL_inst_dft.ap_done == 1'b1)
        region_0_done_cnt <= region_0_done_cnt + 32'h1;
    else;
end


    df_process_intf process_intf_1(clock,reset);
    assign process_intf_1.ap_start = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_start;
    assign process_intf_1.ap_ready = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_ready;
    assign process_intf_1.ap_done = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_done;
    assign process_intf_1.ap_continue = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_continue;
    assign process_intf_1.real_start = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_start;
    assign process_intf_1.pin_stall = 1'b0;
    assign process_intf_1.pout_stall = 1'b0;
    assign process_intf_1.cin_stall = 1'b0;
    assign process_intf_1.cout_stall = 1'b0;
    assign process_intf_1.region_idle = region_0_idle;
    assign process_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_1;
    csv_file_dump pstatus_csv_dumper_1;
    df_process_monitor process_monitor_1;
    df_process_intf process_intf_2(clock,reset);
    assign process_intf_2.ap_start = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_start;
    assign process_intf_2.ap_ready = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_ready;
    assign process_intf_2.ap_done = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_done;
    assign process_intf_2.ap_continue = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_continue;
    assign process_intf_2.real_start = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.ap_start;
    assign process_intf_2.pin_stall = 1'b0;
    assign process_intf_2.pout_stall = 1'b0;
    assign process_intf_2.cin_stall = 1'b0;
    assign process_intf_2.cout_stall = 1'b0;
    assign process_intf_2.region_idle = region_0_idle;
    assign process_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_2;
    csv_file_dump pstatus_csv_dumper_2;
    df_process_monitor process_monitor_2;

    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_dft.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_dft.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_dft.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;

    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.quit_enable = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.loop_start = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_done;
    assign upc_loop_intf_1.loop_continue = AESL_inst_dft.Loop_VITIS_LOOP_16_1_proc_U0.ap_continue;
    assign upc_loop_intf_1.quit_at_end = 1'b0;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.quit_state = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_enable_reg_pp0_iter1282;
    assign upc_loop_intf_2.quit_enable = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_enable_reg_pp0_iter1282;
    assign upc_loop_intf_2.loop_start = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_dft.Loop_VITIS_LOOP_21_2_proc_U0.grp_Loop_VITIS_LOOP_21_2_proc_Pipeline_VITIS_LOOP_21_2_fu_2072.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(1) upc_loop_monitor_2;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;

    fifo_csv_dumper_1 = new("./depth1.csv");
    cstatus_csv_dumper_1 = new("./chan_status1.csv");
    fifo_monitor_1 = new(fifo_csv_dumper_1,fifo_intf_1,cstatus_csv_dumper_1);
    fifo_csv_dumper_2 = new("./depth2.csv");
    cstatus_csv_dumper_2 = new("./chan_status2.csv");
    fifo_monitor_2 = new(fifo_csv_dumper_2,fifo_intf_2,cstatus_csv_dumper_2);
    fifo_csv_dumper_3 = new("./depth3.csv");
    cstatus_csv_dumper_3 = new("./chan_status3.csv");
    fifo_monitor_3 = new(fifo_csv_dumper_3,fifo_intf_3,cstatus_csv_dumper_3);
    fifo_csv_dumper_4 = new("./depth4.csv");
    cstatus_csv_dumper_4 = new("./chan_status4.csv");
    fifo_monitor_4 = new(fifo_csv_dumper_4,fifo_intf_4,cstatus_csv_dumper_4);
    fifo_csv_dumper_5 = new("./depth5.csv");
    cstatus_csv_dumper_5 = new("./chan_status5.csv");
    fifo_monitor_5 = new(fifo_csv_dumper_5,fifo_intf_5,cstatus_csv_dumper_5);
    fifo_csv_dumper_6 = new("./depth6.csv");
    cstatus_csv_dumper_6 = new("./chan_status6.csv");
    fifo_monitor_6 = new(fifo_csv_dumper_6,fifo_intf_6,cstatus_csv_dumper_6);
    fifo_csv_dumper_7 = new("./depth7.csv");
    cstatus_csv_dumper_7 = new("./chan_status7.csv");
    fifo_monitor_7 = new(fifo_csv_dumper_7,fifo_intf_7,cstatus_csv_dumper_7);
    fifo_csv_dumper_8 = new("./depth8.csv");
    cstatus_csv_dumper_8 = new("./chan_status8.csv");
    fifo_monitor_8 = new(fifo_csv_dumper_8,fifo_intf_8,cstatus_csv_dumper_8);
    fifo_csv_dumper_9 = new("./depth9.csv");
    cstatus_csv_dumper_9 = new("./chan_status9.csv");
    fifo_monitor_9 = new(fifo_csv_dumper_9,fifo_intf_9,cstatus_csv_dumper_9);
    fifo_csv_dumper_10 = new("./depth10.csv");
    cstatus_csv_dumper_10 = new("./chan_status10.csv");
    fifo_monitor_10 = new(fifo_csv_dumper_10,fifo_intf_10,cstatus_csv_dumper_10);
    fifo_csv_dumper_11 = new("./depth11.csv");
    cstatus_csv_dumper_11 = new("./chan_status11.csv");
    fifo_monitor_11 = new(fifo_csv_dumper_11,fifo_intf_11,cstatus_csv_dumper_11);
    fifo_csv_dumper_12 = new("./depth12.csv");
    cstatus_csv_dumper_12 = new("./chan_status12.csv");
    fifo_monitor_12 = new(fifo_csv_dumper_12,fifo_intf_12,cstatus_csv_dumper_12);
    fifo_csv_dumper_13 = new("./depth13.csv");
    cstatus_csv_dumper_13 = new("./chan_status13.csv");
    fifo_monitor_13 = new(fifo_csv_dumper_13,fifo_intf_13,cstatus_csv_dumper_13);
    fifo_csv_dumper_14 = new("./depth14.csv");
    cstatus_csv_dumper_14 = new("./chan_status14.csv");
    fifo_monitor_14 = new(fifo_csv_dumper_14,fifo_intf_14,cstatus_csv_dumper_14);
    fifo_csv_dumper_15 = new("./depth15.csv");
    cstatus_csv_dumper_15 = new("./chan_status15.csv");
    fifo_monitor_15 = new(fifo_csv_dumper_15,fifo_intf_15,cstatus_csv_dumper_15);
    fifo_csv_dumper_16 = new("./depth16.csv");
    cstatus_csv_dumper_16 = new("./chan_status16.csv");
    fifo_monitor_16 = new(fifo_csv_dumper_16,fifo_intf_16,cstatus_csv_dumper_16);
    fifo_csv_dumper_17 = new("./depth17.csv");
    cstatus_csv_dumper_17 = new("./chan_status17.csv");
    fifo_monitor_17 = new(fifo_csv_dumper_17,fifo_intf_17,cstatus_csv_dumper_17);
    fifo_csv_dumper_18 = new("./depth18.csv");
    cstatus_csv_dumper_18 = new("./chan_status18.csv");
    fifo_monitor_18 = new(fifo_csv_dumper_18,fifo_intf_18,cstatus_csv_dumper_18);
    fifo_csv_dumper_19 = new("./depth19.csv");
    cstatus_csv_dumper_19 = new("./chan_status19.csv");
    fifo_monitor_19 = new(fifo_csv_dumper_19,fifo_intf_19,cstatus_csv_dumper_19);
    fifo_csv_dumper_20 = new("./depth20.csv");
    cstatus_csv_dumper_20 = new("./chan_status20.csv");
    fifo_monitor_20 = new(fifo_csv_dumper_20,fifo_intf_20,cstatus_csv_dumper_20);
    fifo_csv_dumper_21 = new("./depth21.csv");
    cstatus_csv_dumper_21 = new("./chan_status21.csv");
    fifo_monitor_21 = new(fifo_csv_dumper_21,fifo_intf_21,cstatus_csv_dumper_21);
    fifo_csv_dumper_22 = new("./depth22.csv");
    cstatus_csv_dumper_22 = new("./chan_status22.csv");
    fifo_monitor_22 = new(fifo_csv_dumper_22,fifo_intf_22,cstatus_csv_dumper_22);
    fifo_csv_dumper_23 = new("./depth23.csv");
    cstatus_csv_dumper_23 = new("./chan_status23.csv");
    fifo_monitor_23 = new(fifo_csv_dumper_23,fifo_intf_23,cstatus_csv_dumper_23);
    fifo_csv_dumper_24 = new("./depth24.csv");
    cstatus_csv_dumper_24 = new("./chan_status24.csv");
    fifo_monitor_24 = new(fifo_csv_dumper_24,fifo_intf_24,cstatus_csv_dumper_24);
    fifo_csv_dumper_25 = new("./depth25.csv");
    cstatus_csv_dumper_25 = new("./chan_status25.csv");
    fifo_monitor_25 = new(fifo_csv_dumper_25,fifo_intf_25,cstatus_csv_dumper_25);
    fifo_csv_dumper_26 = new("./depth26.csv");
    cstatus_csv_dumper_26 = new("./chan_status26.csv");
    fifo_monitor_26 = new(fifo_csv_dumper_26,fifo_intf_26,cstatus_csv_dumper_26);
    fifo_csv_dumper_27 = new("./depth27.csv");
    cstatus_csv_dumper_27 = new("./chan_status27.csv");
    fifo_monitor_27 = new(fifo_csv_dumper_27,fifo_intf_27,cstatus_csv_dumper_27);
    fifo_csv_dumper_28 = new("./depth28.csv");
    cstatus_csv_dumper_28 = new("./chan_status28.csv");
    fifo_monitor_28 = new(fifo_csv_dumper_28,fifo_intf_28,cstatus_csv_dumper_28);
    fifo_csv_dumper_29 = new("./depth29.csv");
    cstatus_csv_dumper_29 = new("./chan_status29.csv");
    fifo_monitor_29 = new(fifo_csv_dumper_29,fifo_intf_29,cstatus_csv_dumper_29);
    fifo_csv_dumper_30 = new("./depth30.csv");
    cstatus_csv_dumper_30 = new("./chan_status30.csv");
    fifo_monitor_30 = new(fifo_csv_dumper_30,fifo_intf_30,cstatus_csv_dumper_30);
    fifo_csv_dumper_31 = new("./depth31.csv");
    cstatus_csv_dumper_31 = new("./chan_status31.csv");
    fifo_monitor_31 = new(fifo_csv_dumper_31,fifo_intf_31,cstatus_csv_dumper_31);
    fifo_csv_dumper_32 = new("./depth32.csv");
    cstatus_csv_dumper_32 = new("./chan_status32.csv");
    fifo_monitor_32 = new(fifo_csv_dumper_32,fifo_intf_32,cstatus_csv_dumper_32);
    fifo_csv_dumper_33 = new("./depth33.csv");
    cstatus_csv_dumper_33 = new("./chan_status33.csv");
    fifo_monitor_33 = new(fifo_csv_dumper_33,fifo_intf_33,cstatus_csv_dumper_33);
    fifo_csv_dumper_34 = new("./depth34.csv");
    cstatus_csv_dumper_34 = new("./chan_status34.csv");
    fifo_monitor_34 = new(fifo_csv_dumper_34,fifo_intf_34,cstatus_csv_dumper_34);
    fifo_csv_dumper_35 = new("./depth35.csv");
    cstatus_csv_dumper_35 = new("./chan_status35.csv");
    fifo_monitor_35 = new(fifo_csv_dumper_35,fifo_intf_35,cstatus_csv_dumper_35);
    fifo_csv_dumper_36 = new("./depth36.csv");
    cstatus_csv_dumper_36 = new("./chan_status36.csv");
    fifo_monitor_36 = new(fifo_csv_dumper_36,fifo_intf_36,cstatus_csv_dumper_36);
    fifo_csv_dumper_37 = new("./depth37.csv");
    cstatus_csv_dumper_37 = new("./chan_status37.csv");
    fifo_monitor_37 = new(fifo_csv_dumper_37,fifo_intf_37,cstatus_csv_dumper_37);
    fifo_csv_dumper_38 = new("./depth38.csv");
    cstatus_csv_dumper_38 = new("./chan_status38.csv");
    fifo_monitor_38 = new(fifo_csv_dumper_38,fifo_intf_38,cstatus_csv_dumper_38);
    fifo_csv_dumper_39 = new("./depth39.csv");
    cstatus_csv_dumper_39 = new("./chan_status39.csv");
    fifo_monitor_39 = new(fifo_csv_dumper_39,fifo_intf_39,cstatus_csv_dumper_39);
    fifo_csv_dumper_40 = new("./depth40.csv");
    cstatus_csv_dumper_40 = new("./chan_status40.csv");
    fifo_monitor_40 = new(fifo_csv_dumper_40,fifo_intf_40,cstatus_csv_dumper_40);
    fifo_csv_dumper_41 = new("./depth41.csv");
    cstatus_csv_dumper_41 = new("./chan_status41.csv");
    fifo_monitor_41 = new(fifo_csv_dumper_41,fifo_intf_41,cstatus_csv_dumper_41);
    fifo_csv_dumper_42 = new("./depth42.csv");
    cstatus_csv_dumper_42 = new("./chan_status42.csv");
    fifo_monitor_42 = new(fifo_csv_dumper_42,fifo_intf_42,cstatus_csv_dumper_42);
    fifo_csv_dumper_43 = new("./depth43.csv");
    cstatus_csv_dumper_43 = new("./chan_status43.csv");
    fifo_monitor_43 = new(fifo_csv_dumper_43,fifo_intf_43,cstatus_csv_dumper_43);
    fifo_csv_dumper_44 = new("./depth44.csv");
    cstatus_csv_dumper_44 = new("./chan_status44.csv");
    fifo_monitor_44 = new(fifo_csv_dumper_44,fifo_intf_44,cstatus_csv_dumper_44);
    fifo_csv_dumper_45 = new("./depth45.csv");
    cstatus_csv_dumper_45 = new("./chan_status45.csv");
    fifo_monitor_45 = new(fifo_csv_dumper_45,fifo_intf_45,cstatus_csv_dumper_45);
    fifo_csv_dumper_46 = new("./depth46.csv");
    cstatus_csv_dumper_46 = new("./chan_status46.csv");
    fifo_monitor_46 = new(fifo_csv_dumper_46,fifo_intf_46,cstatus_csv_dumper_46);
    fifo_csv_dumper_47 = new("./depth47.csv");
    cstatus_csv_dumper_47 = new("./chan_status47.csv");
    fifo_monitor_47 = new(fifo_csv_dumper_47,fifo_intf_47,cstatus_csv_dumper_47);
    fifo_csv_dumper_48 = new("./depth48.csv");
    cstatus_csv_dumper_48 = new("./chan_status48.csv");
    fifo_monitor_48 = new(fifo_csv_dumper_48,fifo_intf_48,cstatus_csv_dumper_48);
    fifo_csv_dumper_49 = new("./depth49.csv");
    cstatus_csv_dumper_49 = new("./chan_status49.csv");
    fifo_monitor_49 = new(fifo_csv_dumper_49,fifo_intf_49,cstatus_csv_dumper_49);
    fifo_csv_dumper_50 = new("./depth50.csv");
    cstatus_csv_dumper_50 = new("./chan_status50.csv");
    fifo_monitor_50 = new(fifo_csv_dumper_50,fifo_intf_50,cstatus_csv_dumper_50);
    fifo_csv_dumper_51 = new("./depth51.csv");
    cstatus_csv_dumper_51 = new("./chan_status51.csv");
    fifo_monitor_51 = new(fifo_csv_dumper_51,fifo_intf_51,cstatus_csv_dumper_51);
    fifo_csv_dumper_52 = new("./depth52.csv");
    cstatus_csv_dumper_52 = new("./chan_status52.csv");
    fifo_monitor_52 = new(fifo_csv_dumper_52,fifo_intf_52,cstatus_csv_dumper_52);
    fifo_csv_dumper_53 = new("./depth53.csv");
    cstatus_csv_dumper_53 = new("./chan_status53.csv");
    fifo_monitor_53 = new(fifo_csv_dumper_53,fifo_intf_53,cstatus_csv_dumper_53);
    fifo_csv_dumper_54 = new("./depth54.csv");
    cstatus_csv_dumper_54 = new("./chan_status54.csv");
    fifo_monitor_54 = new(fifo_csv_dumper_54,fifo_intf_54,cstatus_csv_dumper_54);
    fifo_csv_dumper_55 = new("./depth55.csv");
    cstatus_csv_dumper_55 = new("./chan_status55.csv");
    fifo_monitor_55 = new(fifo_csv_dumper_55,fifo_intf_55,cstatus_csv_dumper_55);
    fifo_csv_dumper_56 = new("./depth56.csv");
    cstatus_csv_dumper_56 = new("./chan_status56.csv");
    fifo_monitor_56 = new(fifo_csv_dumper_56,fifo_intf_56,cstatus_csv_dumper_56);
    fifo_csv_dumper_57 = new("./depth57.csv");
    cstatus_csv_dumper_57 = new("./chan_status57.csv");
    fifo_monitor_57 = new(fifo_csv_dumper_57,fifo_intf_57,cstatus_csv_dumper_57);
    fifo_csv_dumper_58 = new("./depth58.csv");
    cstatus_csv_dumper_58 = new("./chan_status58.csv");
    fifo_monitor_58 = new(fifo_csv_dumper_58,fifo_intf_58,cstatus_csv_dumper_58);
    fifo_csv_dumper_59 = new("./depth59.csv");
    cstatus_csv_dumper_59 = new("./chan_status59.csv");
    fifo_monitor_59 = new(fifo_csv_dumper_59,fifo_intf_59,cstatus_csv_dumper_59);
    fifo_csv_dumper_60 = new("./depth60.csv");
    cstatus_csv_dumper_60 = new("./chan_status60.csv");
    fifo_monitor_60 = new(fifo_csv_dumper_60,fifo_intf_60,cstatus_csv_dumper_60);
    fifo_csv_dumper_61 = new("./depth61.csv");
    cstatus_csv_dumper_61 = new("./chan_status61.csv");
    fifo_monitor_61 = new(fifo_csv_dumper_61,fifo_intf_61,cstatus_csv_dumper_61);
    fifo_csv_dumper_62 = new("./depth62.csv");
    cstatus_csv_dumper_62 = new("./chan_status62.csv");
    fifo_monitor_62 = new(fifo_csv_dumper_62,fifo_intf_62,cstatus_csv_dumper_62);
    fifo_csv_dumper_63 = new("./depth63.csv");
    cstatus_csv_dumper_63 = new("./chan_status63.csv");
    fifo_monitor_63 = new(fifo_csv_dumper_63,fifo_intf_63,cstatus_csv_dumper_63);
    fifo_csv_dumper_64 = new("./depth64.csv");
    cstatus_csv_dumper_64 = new("./chan_status64.csv");
    fifo_monitor_64 = new(fifo_csv_dumper_64,fifo_intf_64,cstatus_csv_dumper_64);
    fifo_csv_dumper_65 = new("./depth65.csv");
    cstatus_csv_dumper_65 = new("./chan_status65.csv");
    fifo_monitor_65 = new(fifo_csv_dumper_65,fifo_intf_65,cstatus_csv_dumper_65);
    fifo_csv_dumper_66 = new("./depth66.csv");
    cstatus_csv_dumper_66 = new("./chan_status66.csv");
    fifo_monitor_66 = new(fifo_csv_dumper_66,fifo_intf_66,cstatus_csv_dumper_66);
    fifo_csv_dumper_67 = new("./depth67.csv");
    cstatus_csv_dumper_67 = new("./chan_status67.csv");
    fifo_monitor_67 = new(fifo_csv_dumper_67,fifo_intf_67,cstatus_csv_dumper_67);
    fifo_csv_dumper_68 = new("./depth68.csv");
    cstatus_csv_dumper_68 = new("./chan_status68.csv");
    fifo_monitor_68 = new(fifo_csv_dumper_68,fifo_intf_68,cstatus_csv_dumper_68);
    fifo_csv_dumper_69 = new("./depth69.csv");
    cstatus_csv_dumper_69 = new("./chan_status69.csv");
    fifo_monitor_69 = new(fifo_csv_dumper_69,fifo_intf_69,cstatus_csv_dumper_69);
    fifo_csv_dumper_70 = new("./depth70.csv");
    cstatus_csv_dumper_70 = new("./chan_status70.csv");
    fifo_monitor_70 = new(fifo_csv_dumper_70,fifo_intf_70,cstatus_csv_dumper_70);
    fifo_csv_dumper_71 = new("./depth71.csv");
    cstatus_csv_dumper_71 = new("./chan_status71.csv");
    fifo_monitor_71 = new(fifo_csv_dumper_71,fifo_intf_71,cstatus_csv_dumper_71);
    fifo_csv_dumper_72 = new("./depth72.csv");
    cstatus_csv_dumper_72 = new("./chan_status72.csv");
    fifo_monitor_72 = new(fifo_csv_dumper_72,fifo_intf_72,cstatus_csv_dumper_72);
    fifo_csv_dumper_73 = new("./depth73.csv");
    cstatus_csv_dumper_73 = new("./chan_status73.csv");
    fifo_monitor_73 = new(fifo_csv_dumper_73,fifo_intf_73,cstatus_csv_dumper_73);
    fifo_csv_dumper_74 = new("./depth74.csv");
    cstatus_csv_dumper_74 = new("./chan_status74.csv");
    fifo_monitor_74 = new(fifo_csv_dumper_74,fifo_intf_74,cstatus_csv_dumper_74);
    fifo_csv_dumper_75 = new("./depth75.csv");
    cstatus_csv_dumper_75 = new("./chan_status75.csv");
    fifo_monitor_75 = new(fifo_csv_dumper_75,fifo_intf_75,cstatus_csv_dumper_75);
    fifo_csv_dumper_76 = new("./depth76.csv");
    cstatus_csv_dumper_76 = new("./chan_status76.csv");
    fifo_monitor_76 = new(fifo_csv_dumper_76,fifo_intf_76,cstatus_csv_dumper_76);
    fifo_csv_dumper_77 = new("./depth77.csv");
    cstatus_csv_dumper_77 = new("./chan_status77.csv");
    fifo_monitor_77 = new(fifo_csv_dumper_77,fifo_intf_77,cstatus_csv_dumper_77);
    fifo_csv_dumper_78 = new("./depth78.csv");
    cstatus_csv_dumper_78 = new("./chan_status78.csv");
    fifo_monitor_78 = new(fifo_csv_dumper_78,fifo_intf_78,cstatus_csv_dumper_78);
    fifo_csv_dumper_79 = new("./depth79.csv");
    cstatus_csv_dumper_79 = new("./chan_status79.csv");
    fifo_monitor_79 = new(fifo_csv_dumper_79,fifo_intf_79,cstatus_csv_dumper_79);
    fifo_csv_dumper_80 = new("./depth80.csv");
    cstatus_csv_dumper_80 = new("./chan_status80.csv");
    fifo_monitor_80 = new(fifo_csv_dumper_80,fifo_intf_80,cstatus_csv_dumper_80);
    fifo_csv_dumper_81 = new("./depth81.csv");
    cstatus_csv_dumper_81 = new("./chan_status81.csv");
    fifo_monitor_81 = new(fifo_csv_dumper_81,fifo_intf_81,cstatus_csv_dumper_81);
    fifo_csv_dumper_82 = new("./depth82.csv");
    cstatus_csv_dumper_82 = new("./chan_status82.csv");
    fifo_monitor_82 = new(fifo_csv_dumper_82,fifo_intf_82,cstatus_csv_dumper_82);
    fifo_csv_dumper_83 = new("./depth83.csv");
    cstatus_csv_dumper_83 = new("./chan_status83.csv");
    fifo_monitor_83 = new(fifo_csv_dumper_83,fifo_intf_83,cstatus_csv_dumper_83);
    fifo_csv_dumper_84 = new("./depth84.csv");
    cstatus_csv_dumper_84 = new("./chan_status84.csv");
    fifo_monitor_84 = new(fifo_csv_dumper_84,fifo_intf_84,cstatus_csv_dumper_84);
    fifo_csv_dumper_85 = new("./depth85.csv");
    cstatus_csv_dumper_85 = new("./chan_status85.csv");
    fifo_monitor_85 = new(fifo_csv_dumper_85,fifo_intf_85,cstatus_csv_dumper_85);
    fifo_csv_dumper_86 = new("./depth86.csv");
    cstatus_csv_dumper_86 = new("./chan_status86.csv");
    fifo_monitor_86 = new(fifo_csv_dumper_86,fifo_intf_86,cstatus_csv_dumper_86);
    fifo_csv_dumper_87 = new("./depth87.csv");
    cstatus_csv_dumper_87 = new("./chan_status87.csv");
    fifo_monitor_87 = new(fifo_csv_dumper_87,fifo_intf_87,cstatus_csv_dumper_87);
    fifo_csv_dumper_88 = new("./depth88.csv");
    cstatus_csv_dumper_88 = new("./chan_status88.csv");
    fifo_monitor_88 = new(fifo_csv_dumper_88,fifo_intf_88,cstatus_csv_dumper_88);
    fifo_csv_dumper_89 = new("./depth89.csv");
    cstatus_csv_dumper_89 = new("./chan_status89.csv");
    fifo_monitor_89 = new(fifo_csv_dumper_89,fifo_intf_89,cstatus_csv_dumper_89);
    fifo_csv_dumper_90 = new("./depth90.csv");
    cstatus_csv_dumper_90 = new("./chan_status90.csv");
    fifo_monitor_90 = new(fifo_csv_dumper_90,fifo_intf_90,cstatus_csv_dumper_90);
    fifo_csv_dumper_91 = new("./depth91.csv");
    cstatus_csv_dumper_91 = new("./chan_status91.csv");
    fifo_monitor_91 = new(fifo_csv_dumper_91,fifo_intf_91,cstatus_csv_dumper_91);
    fifo_csv_dumper_92 = new("./depth92.csv");
    cstatus_csv_dumper_92 = new("./chan_status92.csv");
    fifo_monitor_92 = new(fifo_csv_dumper_92,fifo_intf_92,cstatus_csv_dumper_92);
    fifo_csv_dumper_93 = new("./depth93.csv");
    cstatus_csv_dumper_93 = new("./chan_status93.csv");
    fifo_monitor_93 = new(fifo_csv_dumper_93,fifo_intf_93,cstatus_csv_dumper_93);
    fifo_csv_dumper_94 = new("./depth94.csv");
    cstatus_csv_dumper_94 = new("./chan_status94.csv");
    fifo_monitor_94 = new(fifo_csv_dumper_94,fifo_intf_94,cstatus_csv_dumper_94);
    fifo_csv_dumper_95 = new("./depth95.csv");
    cstatus_csv_dumper_95 = new("./chan_status95.csv");
    fifo_monitor_95 = new(fifo_csv_dumper_95,fifo_intf_95,cstatus_csv_dumper_95);
    fifo_csv_dumper_96 = new("./depth96.csv");
    cstatus_csv_dumper_96 = new("./chan_status96.csv");
    fifo_monitor_96 = new(fifo_csv_dumper_96,fifo_intf_96,cstatus_csv_dumper_96);
    fifo_csv_dumper_97 = new("./depth97.csv");
    cstatus_csv_dumper_97 = new("./chan_status97.csv");
    fifo_monitor_97 = new(fifo_csv_dumper_97,fifo_intf_97,cstatus_csv_dumper_97);
    fifo_csv_dumper_98 = new("./depth98.csv");
    cstatus_csv_dumper_98 = new("./chan_status98.csv");
    fifo_monitor_98 = new(fifo_csv_dumper_98,fifo_intf_98,cstatus_csv_dumper_98);
    fifo_csv_dumper_99 = new("./depth99.csv");
    cstatus_csv_dumper_99 = new("./chan_status99.csv");
    fifo_monitor_99 = new(fifo_csv_dumper_99,fifo_intf_99,cstatus_csv_dumper_99);
    fifo_csv_dumper_100 = new("./depth100.csv");
    cstatus_csv_dumper_100 = new("./chan_status100.csv");
    fifo_monitor_100 = new(fifo_csv_dumper_100,fifo_intf_100,cstatus_csv_dumper_100);
    fifo_csv_dumper_101 = new("./depth101.csv");
    cstatus_csv_dumper_101 = new("./chan_status101.csv");
    fifo_monitor_101 = new(fifo_csv_dumper_101,fifo_intf_101,cstatus_csv_dumper_101);
    fifo_csv_dumper_102 = new("./depth102.csv");
    cstatus_csv_dumper_102 = new("./chan_status102.csv");
    fifo_monitor_102 = new(fifo_csv_dumper_102,fifo_intf_102,cstatus_csv_dumper_102);
    fifo_csv_dumper_103 = new("./depth103.csv");
    cstatus_csv_dumper_103 = new("./chan_status103.csv");
    fifo_monitor_103 = new(fifo_csv_dumper_103,fifo_intf_103,cstatus_csv_dumper_103);
    fifo_csv_dumper_104 = new("./depth104.csv");
    cstatus_csv_dumper_104 = new("./chan_status104.csv");
    fifo_monitor_104 = new(fifo_csv_dumper_104,fifo_intf_104,cstatus_csv_dumper_104);
    fifo_csv_dumper_105 = new("./depth105.csv");
    cstatus_csv_dumper_105 = new("./chan_status105.csv");
    fifo_monitor_105 = new(fifo_csv_dumper_105,fifo_intf_105,cstatus_csv_dumper_105);
    fifo_csv_dumper_106 = new("./depth106.csv");
    cstatus_csv_dumper_106 = new("./chan_status106.csv");
    fifo_monitor_106 = new(fifo_csv_dumper_106,fifo_intf_106,cstatus_csv_dumper_106);
    fifo_csv_dumper_107 = new("./depth107.csv");
    cstatus_csv_dumper_107 = new("./chan_status107.csv");
    fifo_monitor_107 = new(fifo_csv_dumper_107,fifo_intf_107,cstatus_csv_dumper_107);
    fifo_csv_dumper_108 = new("./depth108.csv");
    cstatus_csv_dumper_108 = new("./chan_status108.csv");
    fifo_monitor_108 = new(fifo_csv_dumper_108,fifo_intf_108,cstatus_csv_dumper_108);
    fifo_csv_dumper_109 = new("./depth109.csv");
    cstatus_csv_dumper_109 = new("./chan_status109.csv");
    fifo_monitor_109 = new(fifo_csv_dumper_109,fifo_intf_109,cstatus_csv_dumper_109);
    fifo_csv_dumper_110 = new("./depth110.csv");
    cstatus_csv_dumper_110 = new("./chan_status110.csv");
    fifo_monitor_110 = new(fifo_csv_dumper_110,fifo_intf_110,cstatus_csv_dumper_110);
    fifo_csv_dumper_111 = new("./depth111.csv");
    cstatus_csv_dumper_111 = new("./chan_status111.csv");
    fifo_monitor_111 = new(fifo_csv_dumper_111,fifo_intf_111,cstatus_csv_dumper_111);
    fifo_csv_dumper_112 = new("./depth112.csv");
    cstatus_csv_dumper_112 = new("./chan_status112.csv");
    fifo_monitor_112 = new(fifo_csv_dumper_112,fifo_intf_112,cstatus_csv_dumper_112);
    fifo_csv_dumper_113 = new("./depth113.csv");
    cstatus_csv_dumper_113 = new("./chan_status113.csv");
    fifo_monitor_113 = new(fifo_csv_dumper_113,fifo_intf_113,cstatus_csv_dumper_113);
    fifo_csv_dumper_114 = new("./depth114.csv");
    cstatus_csv_dumper_114 = new("./chan_status114.csv");
    fifo_monitor_114 = new(fifo_csv_dumper_114,fifo_intf_114,cstatus_csv_dumper_114);
    fifo_csv_dumper_115 = new("./depth115.csv");
    cstatus_csv_dumper_115 = new("./chan_status115.csv");
    fifo_monitor_115 = new(fifo_csv_dumper_115,fifo_intf_115,cstatus_csv_dumper_115);
    fifo_csv_dumper_116 = new("./depth116.csv");
    cstatus_csv_dumper_116 = new("./chan_status116.csv");
    fifo_monitor_116 = new(fifo_csv_dumper_116,fifo_intf_116,cstatus_csv_dumper_116);
    fifo_csv_dumper_117 = new("./depth117.csv");
    cstatus_csv_dumper_117 = new("./chan_status117.csv");
    fifo_monitor_117 = new(fifo_csv_dumper_117,fifo_intf_117,cstatus_csv_dumper_117);
    fifo_csv_dumper_118 = new("./depth118.csv");
    cstatus_csv_dumper_118 = new("./chan_status118.csv");
    fifo_monitor_118 = new(fifo_csv_dumper_118,fifo_intf_118,cstatus_csv_dumper_118);
    fifo_csv_dumper_119 = new("./depth119.csv");
    cstatus_csv_dumper_119 = new("./chan_status119.csv");
    fifo_monitor_119 = new(fifo_csv_dumper_119,fifo_intf_119,cstatus_csv_dumper_119);
    fifo_csv_dumper_120 = new("./depth120.csv");
    cstatus_csv_dumper_120 = new("./chan_status120.csv");
    fifo_monitor_120 = new(fifo_csv_dumper_120,fifo_intf_120,cstatus_csv_dumper_120);
    fifo_csv_dumper_121 = new("./depth121.csv");
    cstatus_csv_dumper_121 = new("./chan_status121.csv");
    fifo_monitor_121 = new(fifo_csv_dumper_121,fifo_intf_121,cstatus_csv_dumper_121);
    fifo_csv_dumper_122 = new("./depth122.csv");
    cstatus_csv_dumper_122 = new("./chan_status122.csv");
    fifo_monitor_122 = new(fifo_csv_dumper_122,fifo_intf_122,cstatus_csv_dumper_122);
    fifo_csv_dumper_123 = new("./depth123.csv");
    cstatus_csv_dumper_123 = new("./chan_status123.csv");
    fifo_monitor_123 = new(fifo_csv_dumper_123,fifo_intf_123,cstatus_csv_dumper_123);
    fifo_csv_dumper_124 = new("./depth124.csv");
    cstatus_csv_dumper_124 = new("./chan_status124.csv");
    fifo_monitor_124 = new(fifo_csv_dumper_124,fifo_intf_124,cstatus_csv_dumper_124);
    fifo_csv_dumper_125 = new("./depth125.csv");
    cstatus_csv_dumper_125 = new("./chan_status125.csv");
    fifo_monitor_125 = new(fifo_csv_dumper_125,fifo_intf_125,cstatus_csv_dumper_125);
    fifo_csv_dumper_126 = new("./depth126.csv");
    cstatus_csv_dumper_126 = new("./chan_status126.csv");
    fifo_monitor_126 = new(fifo_csv_dumper_126,fifo_intf_126,cstatus_csv_dumper_126);
    fifo_csv_dumper_127 = new("./depth127.csv");
    cstatus_csv_dumper_127 = new("./chan_status127.csv");
    fifo_monitor_127 = new(fifo_csv_dumper_127,fifo_intf_127,cstatus_csv_dumper_127);
    fifo_csv_dumper_128 = new("./depth128.csv");
    cstatus_csv_dumper_128 = new("./chan_status128.csv");
    fifo_monitor_128 = new(fifo_csv_dumper_128,fifo_intf_128,cstatus_csv_dumper_128);
    fifo_csv_dumper_129 = new("./depth129.csv");
    cstatus_csv_dumper_129 = new("./chan_status129.csv");
    fifo_monitor_129 = new(fifo_csv_dumper_129,fifo_intf_129,cstatus_csv_dumper_129);
    fifo_csv_dumper_130 = new("./depth130.csv");
    cstatus_csv_dumper_130 = new("./chan_status130.csv");
    fifo_monitor_130 = new(fifo_csv_dumper_130,fifo_intf_130,cstatus_csv_dumper_130);
    fifo_csv_dumper_131 = new("./depth131.csv");
    cstatus_csv_dumper_131 = new("./chan_status131.csv");
    fifo_monitor_131 = new(fifo_csv_dumper_131,fifo_intf_131,cstatus_csv_dumper_131);
    fifo_csv_dumper_132 = new("./depth132.csv");
    cstatus_csv_dumper_132 = new("./chan_status132.csv");
    fifo_monitor_132 = new(fifo_csv_dumper_132,fifo_intf_132,cstatus_csv_dumper_132);
    fifo_csv_dumper_133 = new("./depth133.csv");
    cstatus_csv_dumper_133 = new("./chan_status133.csv");
    fifo_monitor_133 = new(fifo_csv_dumper_133,fifo_intf_133,cstatus_csv_dumper_133);
    fifo_csv_dumper_134 = new("./depth134.csv");
    cstatus_csv_dumper_134 = new("./chan_status134.csv");
    fifo_monitor_134 = new(fifo_csv_dumper_134,fifo_intf_134,cstatus_csv_dumper_134);
    fifo_csv_dumper_135 = new("./depth135.csv");
    cstatus_csv_dumper_135 = new("./chan_status135.csv");
    fifo_monitor_135 = new(fifo_csv_dumper_135,fifo_intf_135,cstatus_csv_dumper_135);
    fifo_csv_dumper_136 = new("./depth136.csv");
    cstatus_csv_dumper_136 = new("./chan_status136.csv");
    fifo_monitor_136 = new(fifo_csv_dumper_136,fifo_intf_136,cstatus_csv_dumper_136);
    fifo_csv_dumper_137 = new("./depth137.csv");
    cstatus_csv_dumper_137 = new("./chan_status137.csv");
    fifo_monitor_137 = new(fifo_csv_dumper_137,fifo_intf_137,cstatus_csv_dumper_137);
    fifo_csv_dumper_138 = new("./depth138.csv");
    cstatus_csv_dumper_138 = new("./chan_status138.csv");
    fifo_monitor_138 = new(fifo_csv_dumper_138,fifo_intf_138,cstatus_csv_dumper_138);
    fifo_csv_dumper_139 = new("./depth139.csv");
    cstatus_csv_dumper_139 = new("./chan_status139.csv");
    fifo_monitor_139 = new(fifo_csv_dumper_139,fifo_intf_139,cstatus_csv_dumper_139);
    fifo_csv_dumper_140 = new("./depth140.csv");
    cstatus_csv_dumper_140 = new("./chan_status140.csv");
    fifo_monitor_140 = new(fifo_csv_dumper_140,fifo_intf_140,cstatus_csv_dumper_140);
    fifo_csv_dumper_141 = new("./depth141.csv");
    cstatus_csv_dumper_141 = new("./chan_status141.csv");
    fifo_monitor_141 = new(fifo_csv_dumper_141,fifo_intf_141,cstatus_csv_dumper_141);
    fifo_csv_dumper_142 = new("./depth142.csv");
    cstatus_csv_dumper_142 = new("./chan_status142.csv");
    fifo_monitor_142 = new(fifo_csv_dumper_142,fifo_intf_142,cstatus_csv_dumper_142);
    fifo_csv_dumper_143 = new("./depth143.csv");
    cstatus_csv_dumper_143 = new("./chan_status143.csv");
    fifo_monitor_143 = new(fifo_csv_dumper_143,fifo_intf_143,cstatus_csv_dumper_143);
    fifo_csv_dumper_144 = new("./depth144.csv");
    cstatus_csv_dumper_144 = new("./chan_status144.csv");
    fifo_monitor_144 = new(fifo_csv_dumper_144,fifo_intf_144,cstatus_csv_dumper_144);
    fifo_csv_dumper_145 = new("./depth145.csv");
    cstatus_csv_dumper_145 = new("./chan_status145.csv");
    fifo_monitor_145 = new(fifo_csv_dumper_145,fifo_intf_145,cstatus_csv_dumper_145);
    fifo_csv_dumper_146 = new("./depth146.csv");
    cstatus_csv_dumper_146 = new("./chan_status146.csv");
    fifo_monitor_146 = new(fifo_csv_dumper_146,fifo_intf_146,cstatus_csv_dumper_146);
    fifo_csv_dumper_147 = new("./depth147.csv");
    cstatus_csv_dumper_147 = new("./chan_status147.csv");
    fifo_monitor_147 = new(fifo_csv_dumper_147,fifo_intf_147,cstatus_csv_dumper_147);
    fifo_csv_dumper_148 = new("./depth148.csv");
    cstatus_csv_dumper_148 = new("./chan_status148.csv");
    fifo_monitor_148 = new(fifo_csv_dumper_148,fifo_intf_148,cstatus_csv_dumper_148);
    fifo_csv_dumper_149 = new("./depth149.csv");
    cstatus_csv_dumper_149 = new("./chan_status149.csv");
    fifo_monitor_149 = new(fifo_csv_dumper_149,fifo_intf_149,cstatus_csv_dumper_149);
    fifo_csv_dumper_150 = new("./depth150.csv");
    cstatus_csv_dumper_150 = new("./chan_status150.csv");
    fifo_monitor_150 = new(fifo_csv_dumper_150,fifo_intf_150,cstatus_csv_dumper_150);
    fifo_csv_dumper_151 = new("./depth151.csv");
    cstatus_csv_dumper_151 = new("./chan_status151.csv");
    fifo_monitor_151 = new(fifo_csv_dumper_151,fifo_intf_151,cstatus_csv_dumper_151);
    fifo_csv_dumper_152 = new("./depth152.csv");
    cstatus_csv_dumper_152 = new("./chan_status152.csv");
    fifo_monitor_152 = new(fifo_csv_dumper_152,fifo_intf_152,cstatus_csv_dumper_152);
    fifo_csv_dumper_153 = new("./depth153.csv");
    cstatus_csv_dumper_153 = new("./chan_status153.csv");
    fifo_monitor_153 = new(fifo_csv_dumper_153,fifo_intf_153,cstatus_csv_dumper_153);
    fifo_csv_dumper_154 = new("./depth154.csv");
    cstatus_csv_dumper_154 = new("./chan_status154.csv");
    fifo_monitor_154 = new(fifo_csv_dumper_154,fifo_intf_154,cstatus_csv_dumper_154);
    fifo_csv_dumper_155 = new("./depth155.csv");
    cstatus_csv_dumper_155 = new("./chan_status155.csv");
    fifo_monitor_155 = new(fifo_csv_dumper_155,fifo_intf_155,cstatus_csv_dumper_155);
    fifo_csv_dumper_156 = new("./depth156.csv");
    cstatus_csv_dumper_156 = new("./chan_status156.csv");
    fifo_monitor_156 = new(fifo_csv_dumper_156,fifo_intf_156,cstatus_csv_dumper_156);
    fifo_csv_dumper_157 = new("./depth157.csv");
    cstatus_csv_dumper_157 = new("./chan_status157.csv");
    fifo_monitor_157 = new(fifo_csv_dumper_157,fifo_intf_157,cstatus_csv_dumper_157);
    fifo_csv_dumper_158 = new("./depth158.csv");
    cstatus_csv_dumper_158 = new("./chan_status158.csv");
    fifo_monitor_158 = new(fifo_csv_dumper_158,fifo_intf_158,cstatus_csv_dumper_158);
    fifo_csv_dumper_159 = new("./depth159.csv");
    cstatus_csv_dumper_159 = new("./chan_status159.csv");
    fifo_monitor_159 = new(fifo_csv_dumper_159,fifo_intf_159,cstatus_csv_dumper_159);
    fifo_csv_dumper_160 = new("./depth160.csv");
    cstatus_csv_dumper_160 = new("./chan_status160.csv");
    fifo_monitor_160 = new(fifo_csv_dumper_160,fifo_intf_160,cstatus_csv_dumper_160);
    fifo_csv_dumper_161 = new("./depth161.csv");
    cstatus_csv_dumper_161 = new("./chan_status161.csv");
    fifo_monitor_161 = new(fifo_csv_dumper_161,fifo_intf_161,cstatus_csv_dumper_161);
    fifo_csv_dumper_162 = new("./depth162.csv");
    cstatus_csv_dumper_162 = new("./chan_status162.csv");
    fifo_monitor_162 = new(fifo_csv_dumper_162,fifo_intf_162,cstatus_csv_dumper_162);
    fifo_csv_dumper_163 = new("./depth163.csv");
    cstatus_csv_dumper_163 = new("./chan_status163.csv");
    fifo_monitor_163 = new(fifo_csv_dumper_163,fifo_intf_163,cstatus_csv_dumper_163);
    fifo_csv_dumper_164 = new("./depth164.csv");
    cstatus_csv_dumper_164 = new("./chan_status164.csv");
    fifo_monitor_164 = new(fifo_csv_dumper_164,fifo_intf_164,cstatus_csv_dumper_164);
    fifo_csv_dumper_165 = new("./depth165.csv");
    cstatus_csv_dumper_165 = new("./chan_status165.csv");
    fifo_monitor_165 = new(fifo_csv_dumper_165,fifo_intf_165,cstatus_csv_dumper_165);
    fifo_csv_dumper_166 = new("./depth166.csv");
    cstatus_csv_dumper_166 = new("./chan_status166.csv");
    fifo_monitor_166 = new(fifo_csv_dumper_166,fifo_intf_166,cstatus_csv_dumper_166);
    fifo_csv_dumper_167 = new("./depth167.csv");
    cstatus_csv_dumper_167 = new("./chan_status167.csv");
    fifo_monitor_167 = new(fifo_csv_dumper_167,fifo_intf_167,cstatus_csv_dumper_167);
    fifo_csv_dumper_168 = new("./depth168.csv");
    cstatus_csv_dumper_168 = new("./chan_status168.csv");
    fifo_monitor_168 = new(fifo_csv_dumper_168,fifo_intf_168,cstatus_csv_dumper_168);
    fifo_csv_dumper_169 = new("./depth169.csv");
    cstatus_csv_dumper_169 = new("./chan_status169.csv");
    fifo_monitor_169 = new(fifo_csv_dumper_169,fifo_intf_169,cstatus_csv_dumper_169);
    fifo_csv_dumper_170 = new("./depth170.csv");
    cstatus_csv_dumper_170 = new("./chan_status170.csv");
    fifo_monitor_170 = new(fifo_csv_dumper_170,fifo_intf_170,cstatus_csv_dumper_170);
    fifo_csv_dumper_171 = new("./depth171.csv");
    cstatus_csv_dumper_171 = new("./chan_status171.csv");
    fifo_monitor_171 = new(fifo_csv_dumper_171,fifo_intf_171,cstatus_csv_dumper_171);
    fifo_csv_dumper_172 = new("./depth172.csv");
    cstatus_csv_dumper_172 = new("./chan_status172.csv");
    fifo_monitor_172 = new(fifo_csv_dumper_172,fifo_intf_172,cstatus_csv_dumper_172);
    fifo_csv_dumper_173 = new("./depth173.csv");
    cstatus_csv_dumper_173 = new("./chan_status173.csv");
    fifo_monitor_173 = new(fifo_csv_dumper_173,fifo_intf_173,cstatus_csv_dumper_173);
    fifo_csv_dumper_174 = new("./depth174.csv");
    cstatus_csv_dumper_174 = new("./chan_status174.csv");
    fifo_monitor_174 = new(fifo_csv_dumper_174,fifo_intf_174,cstatus_csv_dumper_174);
    fifo_csv_dumper_175 = new("./depth175.csv");
    cstatus_csv_dumper_175 = new("./chan_status175.csv");
    fifo_monitor_175 = new(fifo_csv_dumper_175,fifo_intf_175,cstatus_csv_dumper_175);
    fifo_csv_dumper_176 = new("./depth176.csv");
    cstatus_csv_dumper_176 = new("./chan_status176.csv");
    fifo_monitor_176 = new(fifo_csv_dumper_176,fifo_intf_176,cstatus_csv_dumper_176);
    fifo_csv_dumper_177 = new("./depth177.csv");
    cstatus_csv_dumper_177 = new("./chan_status177.csv");
    fifo_monitor_177 = new(fifo_csv_dumper_177,fifo_intf_177,cstatus_csv_dumper_177);
    fifo_csv_dumper_178 = new("./depth178.csv");
    cstatus_csv_dumper_178 = new("./chan_status178.csv");
    fifo_monitor_178 = new(fifo_csv_dumper_178,fifo_intf_178,cstatus_csv_dumper_178);
    fifo_csv_dumper_179 = new("./depth179.csv");
    cstatus_csv_dumper_179 = new("./chan_status179.csv");
    fifo_monitor_179 = new(fifo_csv_dumper_179,fifo_intf_179,cstatus_csv_dumper_179);
    fifo_csv_dumper_180 = new("./depth180.csv");
    cstatus_csv_dumper_180 = new("./chan_status180.csv");
    fifo_monitor_180 = new(fifo_csv_dumper_180,fifo_intf_180,cstatus_csv_dumper_180);
    fifo_csv_dumper_181 = new("./depth181.csv");
    cstatus_csv_dumper_181 = new("./chan_status181.csv");
    fifo_monitor_181 = new(fifo_csv_dumper_181,fifo_intf_181,cstatus_csv_dumper_181);
    fifo_csv_dumper_182 = new("./depth182.csv");
    cstatus_csv_dumper_182 = new("./chan_status182.csv");
    fifo_monitor_182 = new(fifo_csv_dumper_182,fifo_intf_182,cstatus_csv_dumper_182);
    fifo_csv_dumper_183 = new("./depth183.csv");
    cstatus_csv_dumper_183 = new("./chan_status183.csv");
    fifo_monitor_183 = new(fifo_csv_dumper_183,fifo_intf_183,cstatus_csv_dumper_183);
    fifo_csv_dumper_184 = new("./depth184.csv");
    cstatus_csv_dumper_184 = new("./chan_status184.csv");
    fifo_monitor_184 = new(fifo_csv_dumper_184,fifo_intf_184,cstatus_csv_dumper_184);
    fifo_csv_dumper_185 = new("./depth185.csv");
    cstatus_csv_dumper_185 = new("./chan_status185.csv");
    fifo_monitor_185 = new(fifo_csv_dumper_185,fifo_intf_185,cstatus_csv_dumper_185);
    fifo_csv_dumper_186 = new("./depth186.csv");
    cstatus_csv_dumper_186 = new("./chan_status186.csv");
    fifo_monitor_186 = new(fifo_csv_dumper_186,fifo_intf_186,cstatus_csv_dumper_186);
    fifo_csv_dumper_187 = new("./depth187.csv");
    cstatus_csv_dumper_187 = new("./chan_status187.csv");
    fifo_monitor_187 = new(fifo_csv_dumper_187,fifo_intf_187,cstatus_csv_dumper_187);
    fifo_csv_dumper_188 = new("./depth188.csv");
    cstatus_csv_dumper_188 = new("./chan_status188.csv");
    fifo_monitor_188 = new(fifo_csv_dumper_188,fifo_intf_188,cstatus_csv_dumper_188);
    fifo_csv_dumper_189 = new("./depth189.csv");
    cstatus_csv_dumper_189 = new("./chan_status189.csv");
    fifo_monitor_189 = new(fifo_csv_dumper_189,fifo_intf_189,cstatus_csv_dumper_189);
    fifo_csv_dumper_190 = new("./depth190.csv");
    cstatus_csv_dumper_190 = new("./chan_status190.csv");
    fifo_monitor_190 = new(fifo_csv_dumper_190,fifo_intf_190,cstatus_csv_dumper_190);
    fifo_csv_dumper_191 = new("./depth191.csv");
    cstatus_csv_dumper_191 = new("./chan_status191.csv");
    fifo_monitor_191 = new(fifo_csv_dumper_191,fifo_intf_191,cstatus_csv_dumper_191);
    fifo_csv_dumper_192 = new("./depth192.csv");
    cstatus_csv_dumper_192 = new("./chan_status192.csv");
    fifo_monitor_192 = new(fifo_csv_dumper_192,fifo_intf_192,cstatus_csv_dumper_192);
    fifo_csv_dumper_193 = new("./depth193.csv");
    cstatus_csv_dumper_193 = new("./chan_status193.csv");
    fifo_monitor_193 = new(fifo_csv_dumper_193,fifo_intf_193,cstatus_csv_dumper_193);
    fifo_csv_dumper_194 = new("./depth194.csv");
    cstatus_csv_dumper_194 = new("./chan_status194.csv");
    fifo_monitor_194 = new(fifo_csv_dumper_194,fifo_intf_194,cstatus_csv_dumper_194);
    fifo_csv_dumper_195 = new("./depth195.csv");
    cstatus_csv_dumper_195 = new("./chan_status195.csv");
    fifo_monitor_195 = new(fifo_csv_dumper_195,fifo_intf_195,cstatus_csv_dumper_195);
    fifo_csv_dumper_196 = new("./depth196.csv");
    cstatus_csv_dumper_196 = new("./chan_status196.csv");
    fifo_monitor_196 = new(fifo_csv_dumper_196,fifo_intf_196,cstatus_csv_dumper_196);
    fifo_csv_dumper_197 = new("./depth197.csv");
    cstatus_csv_dumper_197 = new("./chan_status197.csv");
    fifo_monitor_197 = new(fifo_csv_dumper_197,fifo_intf_197,cstatus_csv_dumper_197);
    fifo_csv_dumper_198 = new("./depth198.csv");
    cstatus_csv_dumper_198 = new("./chan_status198.csv");
    fifo_monitor_198 = new(fifo_csv_dumper_198,fifo_intf_198,cstatus_csv_dumper_198);
    fifo_csv_dumper_199 = new("./depth199.csv");
    cstatus_csv_dumper_199 = new("./chan_status199.csv");
    fifo_monitor_199 = new(fifo_csv_dumper_199,fifo_intf_199,cstatus_csv_dumper_199);
    fifo_csv_dumper_200 = new("./depth200.csv");
    cstatus_csv_dumper_200 = new("./chan_status200.csv");
    fifo_monitor_200 = new(fifo_csv_dumper_200,fifo_intf_200,cstatus_csv_dumper_200);
    fifo_csv_dumper_201 = new("./depth201.csv");
    cstatus_csv_dumper_201 = new("./chan_status201.csv");
    fifo_monitor_201 = new(fifo_csv_dumper_201,fifo_intf_201,cstatus_csv_dumper_201);
    fifo_csv_dumper_202 = new("./depth202.csv");
    cstatus_csv_dumper_202 = new("./chan_status202.csv");
    fifo_monitor_202 = new(fifo_csv_dumper_202,fifo_intf_202,cstatus_csv_dumper_202);
    fifo_csv_dumper_203 = new("./depth203.csv");
    cstatus_csv_dumper_203 = new("./chan_status203.csv");
    fifo_monitor_203 = new(fifo_csv_dumper_203,fifo_intf_203,cstatus_csv_dumper_203);
    fifo_csv_dumper_204 = new("./depth204.csv");
    cstatus_csv_dumper_204 = new("./chan_status204.csv");
    fifo_monitor_204 = new(fifo_csv_dumper_204,fifo_intf_204,cstatus_csv_dumper_204);
    fifo_csv_dumper_205 = new("./depth205.csv");
    cstatus_csv_dumper_205 = new("./chan_status205.csv");
    fifo_monitor_205 = new(fifo_csv_dumper_205,fifo_intf_205,cstatus_csv_dumper_205);
    fifo_csv_dumper_206 = new("./depth206.csv");
    cstatus_csv_dumper_206 = new("./chan_status206.csv");
    fifo_monitor_206 = new(fifo_csv_dumper_206,fifo_intf_206,cstatus_csv_dumper_206);
    fifo_csv_dumper_207 = new("./depth207.csv");
    cstatus_csv_dumper_207 = new("./chan_status207.csv");
    fifo_monitor_207 = new(fifo_csv_dumper_207,fifo_intf_207,cstatus_csv_dumper_207);
    fifo_csv_dumper_208 = new("./depth208.csv");
    cstatus_csv_dumper_208 = new("./chan_status208.csv");
    fifo_monitor_208 = new(fifo_csv_dumper_208,fifo_intf_208,cstatus_csv_dumper_208);
    fifo_csv_dumper_209 = new("./depth209.csv");
    cstatus_csv_dumper_209 = new("./chan_status209.csv");
    fifo_monitor_209 = new(fifo_csv_dumper_209,fifo_intf_209,cstatus_csv_dumper_209);
    fifo_csv_dumper_210 = new("./depth210.csv");
    cstatus_csv_dumper_210 = new("./chan_status210.csv");
    fifo_monitor_210 = new(fifo_csv_dumper_210,fifo_intf_210,cstatus_csv_dumper_210);
    fifo_csv_dumper_211 = new("./depth211.csv");
    cstatus_csv_dumper_211 = new("./chan_status211.csv");
    fifo_monitor_211 = new(fifo_csv_dumper_211,fifo_intf_211,cstatus_csv_dumper_211);
    fifo_csv_dumper_212 = new("./depth212.csv");
    cstatus_csv_dumper_212 = new("./chan_status212.csv");
    fifo_monitor_212 = new(fifo_csv_dumper_212,fifo_intf_212,cstatus_csv_dumper_212);
    fifo_csv_dumper_213 = new("./depth213.csv");
    cstatus_csv_dumper_213 = new("./chan_status213.csv");
    fifo_monitor_213 = new(fifo_csv_dumper_213,fifo_intf_213,cstatus_csv_dumper_213);
    fifo_csv_dumper_214 = new("./depth214.csv");
    cstatus_csv_dumper_214 = new("./chan_status214.csv");
    fifo_monitor_214 = new(fifo_csv_dumper_214,fifo_intf_214,cstatus_csv_dumper_214);
    fifo_csv_dumper_215 = new("./depth215.csv");
    cstatus_csv_dumper_215 = new("./chan_status215.csv");
    fifo_monitor_215 = new(fifo_csv_dumper_215,fifo_intf_215,cstatus_csv_dumper_215);
    fifo_csv_dumper_216 = new("./depth216.csv");
    cstatus_csv_dumper_216 = new("./chan_status216.csv");
    fifo_monitor_216 = new(fifo_csv_dumper_216,fifo_intf_216,cstatus_csv_dumper_216);
    fifo_csv_dumper_217 = new("./depth217.csv");
    cstatus_csv_dumper_217 = new("./chan_status217.csv");
    fifo_monitor_217 = new(fifo_csv_dumper_217,fifo_intf_217,cstatus_csv_dumper_217);
    fifo_csv_dumper_218 = new("./depth218.csv");
    cstatus_csv_dumper_218 = new("./chan_status218.csv");
    fifo_monitor_218 = new(fifo_csv_dumper_218,fifo_intf_218,cstatus_csv_dumper_218);
    fifo_csv_dumper_219 = new("./depth219.csv");
    cstatus_csv_dumper_219 = new("./chan_status219.csv");
    fifo_monitor_219 = new(fifo_csv_dumper_219,fifo_intf_219,cstatus_csv_dumper_219);
    fifo_csv_dumper_220 = new("./depth220.csv");
    cstatus_csv_dumper_220 = new("./chan_status220.csv");
    fifo_monitor_220 = new(fifo_csv_dumper_220,fifo_intf_220,cstatus_csv_dumper_220);
    fifo_csv_dumper_221 = new("./depth221.csv");
    cstatus_csv_dumper_221 = new("./chan_status221.csv");
    fifo_monitor_221 = new(fifo_csv_dumper_221,fifo_intf_221,cstatus_csv_dumper_221);
    fifo_csv_dumper_222 = new("./depth222.csv");
    cstatus_csv_dumper_222 = new("./chan_status222.csv");
    fifo_monitor_222 = new(fifo_csv_dumper_222,fifo_intf_222,cstatus_csv_dumper_222);
    fifo_csv_dumper_223 = new("./depth223.csv");
    cstatus_csv_dumper_223 = new("./chan_status223.csv");
    fifo_monitor_223 = new(fifo_csv_dumper_223,fifo_intf_223,cstatus_csv_dumper_223);
    fifo_csv_dumper_224 = new("./depth224.csv");
    cstatus_csv_dumper_224 = new("./chan_status224.csv");
    fifo_monitor_224 = new(fifo_csv_dumper_224,fifo_intf_224,cstatus_csv_dumper_224);
    fifo_csv_dumper_225 = new("./depth225.csv");
    cstatus_csv_dumper_225 = new("./chan_status225.csv");
    fifo_monitor_225 = new(fifo_csv_dumper_225,fifo_intf_225,cstatus_csv_dumper_225);
    fifo_csv_dumper_226 = new("./depth226.csv");
    cstatus_csv_dumper_226 = new("./chan_status226.csv");
    fifo_monitor_226 = new(fifo_csv_dumper_226,fifo_intf_226,cstatus_csv_dumper_226);
    fifo_csv_dumper_227 = new("./depth227.csv");
    cstatus_csv_dumper_227 = new("./chan_status227.csv");
    fifo_monitor_227 = new(fifo_csv_dumper_227,fifo_intf_227,cstatus_csv_dumper_227);
    fifo_csv_dumper_228 = new("./depth228.csv");
    cstatus_csv_dumper_228 = new("./chan_status228.csv");
    fifo_monitor_228 = new(fifo_csv_dumper_228,fifo_intf_228,cstatus_csv_dumper_228);
    fifo_csv_dumper_229 = new("./depth229.csv");
    cstatus_csv_dumper_229 = new("./chan_status229.csv");
    fifo_monitor_229 = new(fifo_csv_dumper_229,fifo_intf_229,cstatus_csv_dumper_229);
    fifo_csv_dumper_230 = new("./depth230.csv");
    cstatus_csv_dumper_230 = new("./chan_status230.csv");
    fifo_monitor_230 = new(fifo_csv_dumper_230,fifo_intf_230,cstatus_csv_dumper_230);
    fifo_csv_dumper_231 = new("./depth231.csv");
    cstatus_csv_dumper_231 = new("./chan_status231.csv");
    fifo_monitor_231 = new(fifo_csv_dumper_231,fifo_intf_231,cstatus_csv_dumper_231);
    fifo_csv_dumper_232 = new("./depth232.csv");
    cstatus_csv_dumper_232 = new("./chan_status232.csv");
    fifo_monitor_232 = new(fifo_csv_dumper_232,fifo_intf_232,cstatus_csv_dumper_232);
    fifo_csv_dumper_233 = new("./depth233.csv");
    cstatus_csv_dumper_233 = new("./chan_status233.csv");
    fifo_monitor_233 = new(fifo_csv_dumper_233,fifo_intf_233,cstatus_csv_dumper_233);
    fifo_csv_dumper_234 = new("./depth234.csv");
    cstatus_csv_dumper_234 = new("./chan_status234.csv");
    fifo_monitor_234 = new(fifo_csv_dumper_234,fifo_intf_234,cstatus_csv_dumper_234);
    fifo_csv_dumper_235 = new("./depth235.csv");
    cstatus_csv_dumper_235 = new("./chan_status235.csv");
    fifo_monitor_235 = new(fifo_csv_dumper_235,fifo_intf_235,cstatus_csv_dumper_235);
    fifo_csv_dumper_236 = new("./depth236.csv");
    cstatus_csv_dumper_236 = new("./chan_status236.csv");
    fifo_monitor_236 = new(fifo_csv_dumper_236,fifo_intf_236,cstatus_csv_dumper_236);
    fifo_csv_dumper_237 = new("./depth237.csv");
    cstatus_csv_dumper_237 = new("./chan_status237.csv");
    fifo_monitor_237 = new(fifo_csv_dumper_237,fifo_intf_237,cstatus_csv_dumper_237);
    fifo_csv_dumper_238 = new("./depth238.csv");
    cstatus_csv_dumper_238 = new("./chan_status238.csv");
    fifo_monitor_238 = new(fifo_csv_dumper_238,fifo_intf_238,cstatus_csv_dumper_238);
    fifo_csv_dumper_239 = new("./depth239.csv");
    cstatus_csv_dumper_239 = new("./chan_status239.csv");
    fifo_monitor_239 = new(fifo_csv_dumper_239,fifo_intf_239,cstatus_csv_dumper_239);
    fifo_csv_dumper_240 = new("./depth240.csv");
    cstatus_csv_dumper_240 = new("./chan_status240.csv");
    fifo_monitor_240 = new(fifo_csv_dumper_240,fifo_intf_240,cstatus_csv_dumper_240);
    fifo_csv_dumper_241 = new("./depth241.csv");
    cstatus_csv_dumper_241 = new("./chan_status241.csv");
    fifo_monitor_241 = new(fifo_csv_dumper_241,fifo_intf_241,cstatus_csv_dumper_241);
    fifo_csv_dumper_242 = new("./depth242.csv");
    cstatus_csv_dumper_242 = new("./chan_status242.csv");
    fifo_monitor_242 = new(fifo_csv_dumper_242,fifo_intf_242,cstatus_csv_dumper_242);
    fifo_csv_dumper_243 = new("./depth243.csv");
    cstatus_csv_dumper_243 = new("./chan_status243.csv");
    fifo_monitor_243 = new(fifo_csv_dumper_243,fifo_intf_243,cstatus_csv_dumper_243);
    fifo_csv_dumper_244 = new("./depth244.csv");
    cstatus_csv_dumper_244 = new("./chan_status244.csv");
    fifo_monitor_244 = new(fifo_csv_dumper_244,fifo_intf_244,cstatus_csv_dumper_244);
    fifo_csv_dumper_245 = new("./depth245.csv");
    cstatus_csv_dumper_245 = new("./chan_status245.csv");
    fifo_monitor_245 = new(fifo_csv_dumper_245,fifo_intf_245,cstatus_csv_dumper_245);
    fifo_csv_dumper_246 = new("./depth246.csv");
    cstatus_csv_dumper_246 = new("./chan_status246.csv");
    fifo_monitor_246 = new(fifo_csv_dumper_246,fifo_intf_246,cstatus_csv_dumper_246);
    fifo_csv_dumper_247 = new("./depth247.csv");
    cstatus_csv_dumper_247 = new("./chan_status247.csv");
    fifo_monitor_247 = new(fifo_csv_dumper_247,fifo_intf_247,cstatus_csv_dumper_247);
    fifo_csv_dumper_248 = new("./depth248.csv");
    cstatus_csv_dumper_248 = new("./chan_status248.csv");
    fifo_monitor_248 = new(fifo_csv_dumper_248,fifo_intf_248,cstatus_csv_dumper_248);
    fifo_csv_dumper_249 = new("./depth249.csv");
    cstatus_csv_dumper_249 = new("./chan_status249.csv");
    fifo_monitor_249 = new(fifo_csv_dumper_249,fifo_intf_249,cstatus_csv_dumper_249);
    fifo_csv_dumper_250 = new("./depth250.csv");
    cstatus_csv_dumper_250 = new("./chan_status250.csv");
    fifo_monitor_250 = new(fifo_csv_dumper_250,fifo_intf_250,cstatus_csv_dumper_250);
    fifo_csv_dumper_251 = new("./depth251.csv");
    cstatus_csv_dumper_251 = new("./chan_status251.csv");
    fifo_monitor_251 = new(fifo_csv_dumper_251,fifo_intf_251,cstatus_csv_dumper_251);
    fifo_csv_dumper_252 = new("./depth252.csv");
    cstatus_csv_dumper_252 = new("./chan_status252.csv");
    fifo_monitor_252 = new(fifo_csv_dumper_252,fifo_intf_252,cstatus_csv_dumper_252);
    fifo_csv_dumper_253 = new("./depth253.csv");
    cstatus_csv_dumper_253 = new("./chan_status253.csv");
    fifo_monitor_253 = new(fifo_csv_dumper_253,fifo_intf_253,cstatus_csv_dumper_253);
    fifo_csv_dumper_254 = new("./depth254.csv");
    cstatus_csv_dumper_254 = new("./chan_status254.csv");
    fifo_monitor_254 = new(fifo_csv_dumper_254,fifo_intf_254,cstatus_csv_dumper_254);
    fifo_csv_dumper_255 = new("./depth255.csv");
    cstatus_csv_dumper_255 = new("./chan_status255.csv");
    fifo_monitor_255 = new(fifo_csv_dumper_255,fifo_intf_255,cstatus_csv_dumper_255);
    fifo_csv_dumper_256 = new("./depth256.csv");
    cstatus_csv_dumper_256 = new("./chan_status256.csv");
    fifo_monitor_256 = new(fifo_csv_dumper_256,fifo_intf_256,cstatus_csv_dumper_256);

    pstall_csv_dumper_1 = new("./stalling1.csv");
    pstatus_csv_dumper_1 = new("./status1.csv");
    process_monitor_1 = new(pstall_csv_dumper_1,process_intf_1,pstatus_csv_dumper_1);
    pstall_csv_dumper_2 = new("./stalling2.csv");
    pstatus_csv_dumper_2 = new("./status2.csv");
    process_monitor_2 = new(pstall_csv_dumper_2,process_intf_2,pstatus_csv_dumper_2);

    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);




    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);

    sample_manager_inst.add_one_monitor(fifo_monitor_1);
    sample_manager_inst.add_one_monitor(fifo_monitor_2);
    sample_manager_inst.add_one_monitor(fifo_monitor_3);
    sample_manager_inst.add_one_monitor(fifo_monitor_4);
    sample_manager_inst.add_one_monitor(fifo_monitor_5);
    sample_manager_inst.add_one_monitor(fifo_monitor_6);
    sample_manager_inst.add_one_monitor(fifo_monitor_7);
    sample_manager_inst.add_one_monitor(fifo_monitor_8);
    sample_manager_inst.add_one_monitor(fifo_monitor_9);
    sample_manager_inst.add_one_monitor(fifo_monitor_10);
    sample_manager_inst.add_one_monitor(fifo_monitor_11);
    sample_manager_inst.add_one_monitor(fifo_monitor_12);
    sample_manager_inst.add_one_monitor(fifo_monitor_13);
    sample_manager_inst.add_one_monitor(fifo_monitor_14);
    sample_manager_inst.add_one_monitor(fifo_monitor_15);
    sample_manager_inst.add_one_monitor(fifo_monitor_16);
    sample_manager_inst.add_one_monitor(fifo_monitor_17);
    sample_manager_inst.add_one_monitor(fifo_monitor_18);
    sample_manager_inst.add_one_monitor(fifo_monitor_19);
    sample_manager_inst.add_one_monitor(fifo_monitor_20);
    sample_manager_inst.add_one_monitor(fifo_monitor_21);
    sample_manager_inst.add_one_monitor(fifo_monitor_22);
    sample_manager_inst.add_one_monitor(fifo_monitor_23);
    sample_manager_inst.add_one_monitor(fifo_monitor_24);
    sample_manager_inst.add_one_monitor(fifo_monitor_25);
    sample_manager_inst.add_one_monitor(fifo_monitor_26);
    sample_manager_inst.add_one_monitor(fifo_monitor_27);
    sample_manager_inst.add_one_monitor(fifo_monitor_28);
    sample_manager_inst.add_one_monitor(fifo_monitor_29);
    sample_manager_inst.add_one_monitor(fifo_monitor_30);
    sample_manager_inst.add_one_monitor(fifo_monitor_31);
    sample_manager_inst.add_one_monitor(fifo_monitor_32);
    sample_manager_inst.add_one_monitor(fifo_monitor_33);
    sample_manager_inst.add_one_monitor(fifo_monitor_34);
    sample_manager_inst.add_one_monitor(fifo_monitor_35);
    sample_manager_inst.add_one_monitor(fifo_monitor_36);
    sample_manager_inst.add_one_monitor(fifo_monitor_37);
    sample_manager_inst.add_one_monitor(fifo_monitor_38);
    sample_manager_inst.add_one_monitor(fifo_monitor_39);
    sample_manager_inst.add_one_monitor(fifo_monitor_40);
    sample_manager_inst.add_one_monitor(fifo_monitor_41);
    sample_manager_inst.add_one_monitor(fifo_monitor_42);
    sample_manager_inst.add_one_monitor(fifo_monitor_43);
    sample_manager_inst.add_one_monitor(fifo_monitor_44);
    sample_manager_inst.add_one_monitor(fifo_monitor_45);
    sample_manager_inst.add_one_monitor(fifo_monitor_46);
    sample_manager_inst.add_one_monitor(fifo_monitor_47);
    sample_manager_inst.add_one_monitor(fifo_monitor_48);
    sample_manager_inst.add_one_monitor(fifo_monitor_49);
    sample_manager_inst.add_one_monitor(fifo_monitor_50);
    sample_manager_inst.add_one_monitor(fifo_monitor_51);
    sample_manager_inst.add_one_monitor(fifo_monitor_52);
    sample_manager_inst.add_one_monitor(fifo_monitor_53);
    sample_manager_inst.add_one_monitor(fifo_monitor_54);
    sample_manager_inst.add_one_monitor(fifo_monitor_55);
    sample_manager_inst.add_one_monitor(fifo_monitor_56);
    sample_manager_inst.add_one_monitor(fifo_monitor_57);
    sample_manager_inst.add_one_monitor(fifo_monitor_58);
    sample_manager_inst.add_one_monitor(fifo_monitor_59);
    sample_manager_inst.add_one_monitor(fifo_monitor_60);
    sample_manager_inst.add_one_monitor(fifo_monitor_61);
    sample_manager_inst.add_one_monitor(fifo_monitor_62);
    sample_manager_inst.add_one_monitor(fifo_monitor_63);
    sample_manager_inst.add_one_monitor(fifo_monitor_64);
    sample_manager_inst.add_one_monitor(fifo_monitor_65);
    sample_manager_inst.add_one_monitor(fifo_monitor_66);
    sample_manager_inst.add_one_monitor(fifo_monitor_67);
    sample_manager_inst.add_one_monitor(fifo_monitor_68);
    sample_manager_inst.add_one_monitor(fifo_monitor_69);
    sample_manager_inst.add_one_monitor(fifo_monitor_70);
    sample_manager_inst.add_one_monitor(fifo_monitor_71);
    sample_manager_inst.add_one_monitor(fifo_monitor_72);
    sample_manager_inst.add_one_monitor(fifo_monitor_73);
    sample_manager_inst.add_one_monitor(fifo_monitor_74);
    sample_manager_inst.add_one_monitor(fifo_monitor_75);
    sample_manager_inst.add_one_monitor(fifo_monitor_76);
    sample_manager_inst.add_one_monitor(fifo_monitor_77);
    sample_manager_inst.add_one_monitor(fifo_monitor_78);
    sample_manager_inst.add_one_monitor(fifo_monitor_79);
    sample_manager_inst.add_one_monitor(fifo_monitor_80);
    sample_manager_inst.add_one_monitor(fifo_monitor_81);
    sample_manager_inst.add_one_monitor(fifo_monitor_82);
    sample_manager_inst.add_one_monitor(fifo_monitor_83);
    sample_manager_inst.add_one_monitor(fifo_monitor_84);
    sample_manager_inst.add_one_monitor(fifo_monitor_85);
    sample_manager_inst.add_one_monitor(fifo_monitor_86);
    sample_manager_inst.add_one_monitor(fifo_monitor_87);
    sample_manager_inst.add_one_monitor(fifo_monitor_88);
    sample_manager_inst.add_one_monitor(fifo_monitor_89);
    sample_manager_inst.add_one_monitor(fifo_monitor_90);
    sample_manager_inst.add_one_monitor(fifo_monitor_91);
    sample_manager_inst.add_one_monitor(fifo_monitor_92);
    sample_manager_inst.add_one_monitor(fifo_monitor_93);
    sample_manager_inst.add_one_monitor(fifo_monitor_94);
    sample_manager_inst.add_one_monitor(fifo_monitor_95);
    sample_manager_inst.add_one_monitor(fifo_monitor_96);
    sample_manager_inst.add_one_monitor(fifo_monitor_97);
    sample_manager_inst.add_one_monitor(fifo_monitor_98);
    sample_manager_inst.add_one_monitor(fifo_monitor_99);
    sample_manager_inst.add_one_monitor(fifo_monitor_100);
    sample_manager_inst.add_one_monitor(fifo_monitor_101);
    sample_manager_inst.add_one_monitor(fifo_monitor_102);
    sample_manager_inst.add_one_monitor(fifo_monitor_103);
    sample_manager_inst.add_one_monitor(fifo_monitor_104);
    sample_manager_inst.add_one_monitor(fifo_monitor_105);
    sample_manager_inst.add_one_monitor(fifo_monitor_106);
    sample_manager_inst.add_one_monitor(fifo_monitor_107);
    sample_manager_inst.add_one_monitor(fifo_monitor_108);
    sample_manager_inst.add_one_monitor(fifo_monitor_109);
    sample_manager_inst.add_one_monitor(fifo_monitor_110);
    sample_manager_inst.add_one_monitor(fifo_monitor_111);
    sample_manager_inst.add_one_monitor(fifo_monitor_112);
    sample_manager_inst.add_one_monitor(fifo_monitor_113);
    sample_manager_inst.add_one_monitor(fifo_monitor_114);
    sample_manager_inst.add_one_monitor(fifo_monitor_115);
    sample_manager_inst.add_one_monitor(fifo_monitor_116);
    sample_manager_inst.add_one_monitor(fifo_monitor_117);
    sample_manager_inst.add_one_monitor(fifo_monitor_118);
    sample_manager_inst.add_one_monitor(fifo_monitor_119);
    sample_manager_inst.add_one_monitor(fifo_monitor_120);
    sample_manager_inst.add_one_monitor(fifo_monitor_121);
    sample_manager_inst.add_one_monitor(fifo_monitor_122);
    sample_manager_inst.add_one_monitor(fifo_monitor_123);
    sample_manager_inst.add_one_monitor(fifo_monitor_124);
    sample_manager_inst.add_one_monitor(fifo_monitor_125);
    sample_manager_inst.add_one_monitor(fifo_monitor_126);
    sample_manager_inst.add_one_monitor(fifo_monitor_127);
    sample_manager_inst.add_one_monitor(fifo_monitor_128);
    sample_manager_inst.add_one_monitor(fifo_monitor_129);
    sample_manager_inst.add_one_monitor(fifo_monitor_130);
    sample_manager_inst.add_one_monitor(fifo_monitor_131);
    sample_manager_inst.add_one_monitor(fifo_monitor_132);
    sample_manager_inst.add_one_monitor(fifo_monitor_133);
    sample_manager_inst.add_one_monitor(fifo_monitor_134);
    sample_manager_inst.add_one_monitor(fifo_monitor_135);
    sample_manager_inst.add_one_monitor(fifo_monitor_136);
    sample_manager_inst.add_one_monitor(fifo_monitor_137);
    sample_manager_inst.add_one_monitor(fifo_monitor_138);
    sample_manager_inst.add_one_monitor(fifo_monitor_139);
    sample_manager_inst.add_one_monitor(fifo_monitor_140);
    sample_manager_inst.add_one_monitor(fifo_monitor_141);
    sample_manager_inst.add_one_monitor(fifo_monitor_142);
    sample_manager_inst.add_one_monitor(fifo_monitor_143);
    sample_manager_inst.add_one_monitor(fifo_monitor_144);
    sample_manager_inst.add_one_monitor(fifo_monitor_145);
    sample_manager_inst.add_one_monitor(fifo_monitor_146);
    sample_manager_inst.add_one_monitor(fifo_monitor_147);
    sample_manager_inst.add_one_monitor(fifo_monitor_148);
    sample_manager_inst.add_one_monitor(fifo_monitor_149);
    sample_manager_inst.add_one_monitor(fifo_monitor_150);
    sample_manager_inst.add_one_monitor(fifo_monitor_151);
    sample_manager_inst.add_one_monitor(fifo_monitor_152);
    sample_manager_inst.add_one_monitor(fifo_monitor_153);
    sample_manager_inst.add_one_monitor(fifo_monitor_154);
    sample_manager_inst.add_one_monitor(fifo_monitor_155);
    sample_manager_inst.add_one_monitor(fifo_monitor_156);
    sample_manager_inst.add_one_monitor(fifo_monitor_157);
    sample_manager_inst.add_one_monitor(fifo_monitor_158);
    sample_manager_inst.add_one_monitor(fifo_monitor_159);
    sample_manager_inst.add_one_monitor(fifo_monitor_160);
    sample_manager_inst.add_one_monitor(fifo_monitor_161);
    sample_manager_inst.add_one_monitor(fifo_monitor_162);
    sample_manager_inst.add_one_monitor(fifo_monitor_163);
    sample_manager_inst.add_one_monitor(fifo_monitor_164);
    sample_manager_inst.add_one_monitor(fifo_monitor_165);
    sample_manager_inst.add_one_monitor(fifo_monitor_166);
    sample_manager_inst.add_one_monitor(fifo_monitor_167);
    sample_manager_inst.add_one_monitor(fifo_monitor_168);
    sample_manager_inst.add_one_monitor(fifo_monitor_169);
    sample_manager_inst.add_one_monitor(fifo_monitor_170);
    sample_manager_inst.add_one_monitor(fifo_monitor_171);
    sample_manager_inst.add_one_monitor(fifo_monitor_172);
    sample_manager_inst.add_one_monitor(fifo_monitor_173);
    sample_manager_inst.add_one_monitor(fifo_monitor_174);
    sample_manager_inst.add_one_monitor(fifo_monitor_175);
    sample_manager_inst.add_one_monitor(fifo_monitor_176);
    sample_manager_inst.add_one_monitor(fifo_monitor_177);
    sample_manager_inst.add_one_monitor(fifo_monitor_178);
    sample_manager_inst.add_one_monitor(fifo_monitor_179);
    sample_manager_inst.add_one_monitor(fifo_monitor_180);
    sample_manager_inst.add_one_monitor(fifo_monitor_181);
    sample_manager_inst.add_one_monitor(fifo_monitor_182);
    sample_manager_inst.add_one_monitor(fifo_monitor_183);
    sample_manager_inst.add_one_monitor(fifo_monitor_184);
    sample_manager_inst.add_one_monitor(fifo_monitor_185);
    sample_manager_inst.add_one_monitor(fifo_monitor_186);
    sample_manager_inst.add_one_monitor(fifo_monitor_187);
    sample_manager_inst.add_one_monitor(fifo_monitor_188);
    sample_manager_inst.add_one_monitor(fifo_monitor_189);
    sample_manager_inst.add_one_monitor(fifo_monitor_190);
    sample_manager_inst.add_one_monitor(fifo_monitor_191);
    sample_manager_inst.add_one_monitor(fifo_monitor_192);
    sample_manager_inst.add_one_monitor(fifo_monitor_193);
    sample_manager_inst.add_one_monitor(fifo_monitor_194);
    sample_manager_inst.add_one_monitor(fifo_monitor_195);
    sample_manager_inst.add_one_monitor(fifo_monitor_196);
    sample_manager_inst.add_one_monitor(fifo_monitor_197);
    sample_manager_inst.add_one_monitor(fifo_monitor_198);
    sample_manager_inst.add_one_monitor(fifo_monitor_199);
    sample_manager_inst.add_one_monitor(fifo_monitor_200);
    sample_manager_inst.add_one_monitor(fifo_monitor_201);
    sample_manager_inst.add_one_monitor(fifo_monitor_202);
    sample_manager_inst.add_one_monitor(fifo_monitor_203);
    sample_manager_inst.add_one_monitor(fifo_monitor_204);
    sample_manager_inst.add_one_monitor(fifo_monitor_205);
    sample_manager_inst.add_one_monitor(fifo_monitor_206);
    sample_manager_inst.add_one_monitor(fifo_monitor_207);
    sample_manager_inst.add_one_monitor(fifo_monitor_208);
    sample_manager_inst.add_one_monitor(fifo_monitor_209);
    sample_manager_inst.add_one_monitor(fifo_monitor_210);
    sample_manager_inst.add_one_monitor(fifo_monitor_211);
    sample_manager_inst.add_one_monitor(fifo_monitor_212);
    sample_manager_inst.add_one_monitor(fifo_monitor_213);
    sample_manager_inst.add_one_monitor(fifo_monitor_214);
    sample_manager_inst.add_one_monitor(fifo_monitor_215);
    sample_manager_inst.add_one_monitor(fifo_monitor_216);
    sample_manager_inst.add_one_monitor(fifo_monitor_217);
    sample_manager_inst.add_one_monitor(fifo_monitor_218);
    sample_manager_inst.add_one_monitor(fifo_monitor_219);
    sample_manager_inst.add_one_monitor(fifo_monitor_220);
    sample_manager_inst.add_one_monitor(fifo_monitor_221);
    sample_manager_inst.add_one_monitor(fifo_monitor_222);
    sample_manager_inst.add_one_monitor(fifo_monitor_223);
    sample_manager_inst.add_one_monitor(fifo_monitor_224);
    sample_manager_inst.add_one_monitor(fifo_monitor_225);
    sample_manager_inst.add_one_monitor(fifo_monitor_226);
    sample_manager_inst.add_one_monitor(fifo_monitor_227);
    sample_manager_inst.add_one_monitor(fifo_monitor_228);
    sample_manager_inst.add_one_monitor(fifo_monitor_229);
    sample_manager_inst.add_one_monitor(fifo_monitor_230);
    sample_manager_inst.add_one_monitor(fifo_monitor_231);
    sample_manager_inst.add_one_monitor(fifo_monitor_232);
    sample_manager_inst.add_one_monitor(fifo_monitor_233);
    sample_manager_inst.add_one_monitor(fifo_monitor_234);
    sample_manager_inst.add_one_monitor(fifo_monitor_235);
    sample_manager_inst.add_one_monitor(fifo_monitor_236);
    sample_manager_inst.add_one_monitor(fifo_monitor_237);
    sample_manager_inst.add_one_monitor(fifo_monitor_238);
    sample_manager_inst.add_one_monitor(fifo_monitor_239);
    sample_manager_inst.add_one_monitor(fifo_monitor_240);
    sample_manager_inst.add_one_monitor(fifo_monitor_241);
    sample_manager_inst.add_one_monitor(fifo_monitor_242);
    sample_manager_inst.add_one_monitor(fifo_monitor_243);
    sample_manager_inst.add_one_monitor(fifo_monitor_244);
    sample_manager_inst.add_one_monitor(fifo_monitor_245);
    sample_manager_inst.add_one_monitor(fifo_monitor_246);
    sample_manager_inst.add_one_monitor(fifo_monitor_247);
    sample_manager_inst.add_one_monitor(fifo_monitor_248);
    sample_manager_inst.add_one_monitor(fifo_monitor_249);
    sample_manager_inst.add_one_monitor(fifo_monitor_250);
    sample_manager_inst.add_one_monitor(fifo_monitor_251);
    sample_manager_inst.add_one_monitor(fifo_monitor_252);
    sample_manager_inst.add_one_monitor(fifo_monitor_253);
    sample_manager_inst.add_one_monitor(fifo_monitor_254);
    sample_manager_inst.add_one_monitor(fifo_monitor_255);
    sample_manager_inst.add_one_monitor(fifo_monitor_256);
    sample_manager_inst.add_one_monitor(process_monitor_1);
    sample_manager_inst.add_one_monitor(process_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1 || deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
